library verilog;
use verilog.vl_types.all;
entity TOPLEVEL is
    port(
        CAPTURE         : in     vl_logic;
        CLK50           : in     vl_logic;
        MAC_CRSDV       : in     vl_logic;
        MAC_RXD         : in     vl_logic_vector(1 downto 0);
        MAC_RXER        : in     vl_logic;
        MAINXIN         : in     vl_logic;
        MISO            : in     vl_logic;
        MSS_RESET_N     : in     vl_logic;
        UART_0_RXD      : in     vl_logic;
        CS              : out    vl_logic;
        MAC_MDC         : out    vl_logic;
        MAC_TXD         : out    vl_logic_vector(1 downto 0);
        MAC_TXEN        : out    vl_logic;
        Phy_RMII_CLK    : out    vl_logic;
        SCLK            : out    vl_logic;
        UART_0_TXD      : out    vl_logic;
        adcConvComplete : out    vl_logic;
        adcStartCapture : out    vl_logic;
        incp            : out    vl_logic;
        incv            : out    vl_logic;
        inphi           : out    vl_logic;
        led             : out    vl_logic_vector(7 downto 0);
        psram_address   : out    vl_logic_vector(24 downto 0);
        psram_nbyte_en  : out    vl_logic_vector(1 downto 0);
        psram_ncs0      : out    vl_logic;
        psram_ncs1      : out    vl_logic;
        psram_noe0      : out    vl_logic;
        psram_noe1      : out    vl_logic;
        psram_nwe       : out    vl_logic;
        resp            : out    vl_logic;
        resv            : out    vl_logic;
        rs485_de        : out    vl_logic;
        rs485_nre       : out    vl_logic;
        MAC_MDIO        : inout  vl_logic;
        psram_data      : inout  vl_logic_vector(15 downto 0)
    );
end TOPLEVEL;
