library verilog;
use verilog.vl_types.all;
entity BFM_MAIN is
    generic(
        OPMODE          : integer := 0;
        VECTFILE        : string  := "test.vec";
        MAX_INSTRUCTIONS: integer := 16384;
        MAX_STACK       : integer := 1024;
        MAX_MEMTEST     : integer := 65536;
        TPD             : integer := 1;
        DEBUGLEVEL      : integer := -1;
        CON_SPULSE      : integer := 0;
        ARGVALUE0       : integer := 0;
        ARGVALUE1       : integer := 0;
        ARGVALUE2       : integer := 0;
        ARGVALUE3       : integer := 0;
        ARGVALUE4       : integer := 0;
        ARGVALUE5       : integer := 0;
        ARGVALUE6       : integer := 0;
        ARGVALUE7       : integer := 0;
        ARGVALUE8       : integer := 0;
        ARGVALUE9       : integer := 0;
        ARGVALUE10      : integer := 0;
        ARGVALUE11      : integer := 0;
        ARGVALUE12      : integer := 0;
        ARGVALUE13      : integer := 0;
        ARGVALUE14      : integer := 0;
        ARGVALUE15      : integer := 0;
        ARGVALUE16      : integer := 0;
        ARGVALUE17      : integer := 0;
        ARGVALUE18      : integer := 0;
        ARGVALUE19      : integer := 0;
        ARGVALUE20      : integer := 0;
        ARGVALUE21      : integer := 0;
        ARGVALUE22      : integer := 0;
        ARGVALUE23      : integer := 0;
        ARGVALUE24      : integer := 0;
        ARGVALUE25      : integer := 0;
        ARGVALUE26      : integer := 0;
        ARGVALUE27      : integer := 0;
        ARGVALUE28      : integer := 0;
        ARGVALUE29      : integer := 0;
        ARGVALUE30      : integer := 0;
        ARGVALUE31      : integer := 0;
        ARGVALUE32      : integer := 0;
        ARGVALUE33      : integer := 0;
        ARGVALUE34      : integer := 0;
        ARGVALUE35      : integer := 0;
        ARGVALUE36      : integer := 0;
        ARGVALUE37      : integer := 0;
        ARGVALUE38      : integer := 0;
        ARGVALUE39      : integer := 0;
        ARGVALUE40      : integer := 0;
        ARGVALUE41      : integer := 0;
        ARGVALUE42      : integer := 0;
        ARGVALUE43      : integer := 0;
        ARGVALUE44      : integer := 0;
        ARGVALUE45      : integer := 0;
        ARGVALUE46      : integer := 0;
        ARGVALUE47      : integer := 0;
        ARGVALUE48      : integer := 0;
        ARGVALUE49      : integer := 0;
        ARGVALUE50      : integer := 0;
        ARGVALUE51      : integer := 0;
        ARGVALUE52      : integer := 0;
        ARGVALUE53      : integer := 0;
        ARGVALUE54      : integer := 0;
        ARGVALUE55      : integer := 0;
        ARGVALUE56      : integer := 0;
        ARGVALUE57      : integer := 0;
        ARGVALUE58      : integer := 0;
        ARGVALUE59      : integer := 0;
        ARGVALUE60      : integer := 0;
        ARGVALUE61      : integer := 0;
        ARGVALUE62      : integer := 0;
        ARGVALUE63      : integer := 0;
        ARGVALUE64      : integer := 0;
        ARGVALUE65      : integer := 0;
        ARGVALUE66      : integer := 0;
        ARGVALUE67      : integer := 0;
        ARGVALUE68      : integer := 0;
        ARGVALUE69      : integer := 0;
        ARGVALUE70      : integer := 0;
        ARGVALUE71      : integer := 0;
        ARGVALUE72      : integer := 0;
        ARGVALUE73      : integer := 0;
        ARGVALUE74      : integer := 0;
        ARGVALUE75      : integer := 0;
        ARGVALUE76      : integer := 0;
        ARGVALUE77      : integer := 0;
        ARGVALUE78      : integer := 0;
        ARGVALUE79      : integer := 0;
        ARGVALUE80      : integer := 0;
        ARGVALUE81      : integer := 0;
        ARGVALUE82      : integer := 0;
        ARGVALUE83      : integer := 0;
        ARGVALUE84      : integer := 0;
        ARGVALUE85      : integer := 0;
        ARGVALUE86      : integer := 0;
        ARGVALUE87      : integer := 0;
        ARGVALUE88      : integer := 0;
        ARGVALUE89      : integer := 0;
        ARGVALUE90      : integer := 0;
        ARGVALUE91      : integer := 0;
        ARGVALUE92      : integer := 0;
        ARGVALUE93      : integer := 0;
        ARGVALUE94      : integer := 0;
        ARGVALUE95      : integer := 0;
        ARGVALUE96      : integer := 0;
        ARGVALUE97      : integer := 0;
        ARGVALUE98      : integer := 0;
        ARGVALUE99      : integer := 0;
        ZEROLV          : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ZERO256         : vl_logic_vector(255 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TPDns           : vl_notype;
        idle            : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        init            : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        active          : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        done            : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        fill            : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        scan            : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi1)
    );
    port(
        SYSCLK          : in     vl_logic;
        SYSRSTN         : in     vl_logic;
        PCLK            : out    vl_logic;
        HCLK            : out    vl_logic;
        HRESETN         : out    vl_logic;
        HADDR           : out    vl_logic_vector(31 downto 0);
        HBURST          : out    vl_logic_vector(2 downto 0);
        HMASTLOCK       : out    vl_logic;
        HPROT           : out    vl_logic_vector(3 downto 0);
        HSIZE           : out    vl_logic_vector(2 downto 0);
        HTRANS          : out    vl_logic_vector(1 downto 0);
        HWRITE          : out    vl_logic;
        HWDATA          : out    vl_logic_vector(31 downto 0);
        HRDATA          : in     vl_logic_vector(31 downto 0);
        HREADY          : in     vl_logic;
        HRESP           : in     vl_logic;
        HSEL            : out    vl_logic_vector(15 downto 0);
        INTERRUPT       : in     vl_logic_vector(255 downto 0);
        GP_OUT          : out    vl_logic_vector(31 downto 0);
        GP_IN           : in     vl_logic_vector(31 downto 0);
        EXT_WR          : out    vl_logic;
        EXT_RD          : out    vl_logic;
        EXT_ADDR        : out    vl_logic_vector(31 downto 0);
        EXT_DATA        : inout  vl_logic_vector(31 downto 0);
        EXT_WAIT        : in     vl_logic;
        CON_ADDR        : in     vl_logic_vector(15 downto 0);
        CON_DATA        : inout  vl_logic_vector(31 downto 0);
        CON_RD          : in     vl_logic;
        CON_WR          : in     vl_logic;
        CON_BUSY        : out    vl_logic;
        INSTR_OUT       : out    vl_logic_vector(31 downto 0);
        INSTR_IN        : in     vl_logic_vector(31 downto 0);
        FINISHED        : out    vl_logic;
        FAILED          : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of OPMODE : constant is 1;
    attribute mti_svvh_generic_type of VECTFILE : constant is 1;
    attribute mti_svvh_generic_type of MAX_INSTRUCTIONS : constant is 1;
    attribute mti_svvh_generic_type of MAX_STACK : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEMTEST : constant is 1;
    attribute mti_svvh_generic_type of TPD : constant is 1;
    attribute mti_svvh_generic_type of DEBUGLEVEL : constant is 1;
    attribute mti_svvh_generic_type of CON_SPULSE : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE0 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE1 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE2 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE3 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE4 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE5 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE6 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE7 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE8 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE9 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE10 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE11 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE12 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE13 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE14 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE15 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE16 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE17 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE18 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE19 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE20 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE21 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE22 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE23 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE24 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE25 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE26 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE27 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE28 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE29 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE30 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE31 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE32 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE33 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE34 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE35 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE36 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE37 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE38 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE39 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE40 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE41 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE42 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE43 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE44 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE45 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE46 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE47 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE48 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE49 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE50 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE51 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE52 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE53 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE54 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE55 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE56 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE57 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE58 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE59 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE60 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE61 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE62 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE63 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE64 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE65 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE66 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE67 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE68 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE69 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE70 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE71 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE72 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE73 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE74 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE75 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE76 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE77 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE78 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE79 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE80 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE81 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE82 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE83 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE84 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE85 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE86 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE87 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE88 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE89 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE90 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE91 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE92 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE93 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE94 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE95 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE96 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE97 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE98 : constant is 1;
    attribute mti_svvh_generic_type of ARGVALUE99 : constant is 1;
    attribute mti_svvh_generic_type of ZEROLV : constant is 2;
    attribute mti_svvh_generic_type of ZERO256 : constant is 2;
    attribute mti_svvh_generic_type of TPDns : constant is 3;
    attribute mti_svvh_generic_type of idle : constant is 2;
    attribute mti_svvh_generic_type of init : constant is 2;
    attribute mti_svvh_generic_type of active : constant is 2;
    attribute mti_svvh_generic_type of done : constant is 2;
    attribute mti_svvh_generic_type of fill : constant is 2;
    attribute mti_svvh_generic_type of scan : constant is 2;
end BFM_MAIN;
