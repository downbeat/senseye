library verilog;
use verilog.vl_types.all;
entity F2AB is
    generic(
        WIDTH           : integer := 32;
        DAC_RESOLUTION  : integer := 0;
        WARNING_MSGS_ON : integer := 1;
        FAST_ADC_CONV_SIM: integer := 0;
        ANALOG_QUAD_NUM : integer := 6;
        ADC_NUM         : integer := 3;
        NUM_ADC_IN      : integer := 5;
        VAREF_INT       : real    := 2.560000
    );
    port(
        AV1             : in     vl_logic_vector(5 downto 0);
        AV2             : in     vl_logic_vector(5 downto 0);
        AC              : in     vl_logic_vector(5 downto 0);
        AT              : in     vl_logic_vector(5 downto 0);
        ATGND_01        : in     vl_logic;
        ATGND_23        : in     vl_logic;
        ATGND_45        : in     vl_logic;
        VAREF           : in     vl_logic_vector(2 downto 0);
        ADCGNDREF       : in     vl_logic;
        ADC_VAREFSEL    : in     vl_logic;
        ADC0            : in     vl_logic_vector(3 downto 0);
        ADC1            : in     vl_logic_vector(3 downto 0);
        ADC2            : in     vl_logic_vector(3 downto 0);
        DEN_ADC         : in     vl_logic_vector(11 downto 0);
        ADC0_PWRDWN     : in     vl_logic;
        ADC0_ADCRESET   : in     vl_logic;
        ADC0_SYSCLK     : in     vl_logic;
        ADC0_CHNUMBER   : in     vl_logic_vector(4 downto 0);
        ADC0_MODE       : in     vl_logic_vector(3 downto 0);
        ADC0_TVC        : in     vl_logic_vector(7 downto 0);
        ADC0_STC        : in     vl_logic_vector(7 downto 0);
        ADC0_ADCSTART   : in     vl_logic;
        ADC1_PWRDWN     : in     vl_logic;
        ADC1_ADCRESET   : in     vl_logic;
        ADC1_SYSCLK     : in     vl_logic;
        ADC1_CHNUMBER   : in     vl_logic_vector(4 downto 0);
        ADC1_MODE       : in     vl_logic_vector(3 downto 0);
        ADC1_TVC        : in     vl_logic_vector(7 downto 0);
        ADC1_STC        : in     vl_logic_vector(7 downto 0);
        ADC1_ADCSTART   : in     vl_logic;
        ADC2_PWRDWN     : in     vl_logic;
        ADC2_ADCRESET   : in     vl_logic;
        ADC2_SYSCLK     : in     vl_logic;
        ADC2_CHNUMBER   : in     vl_logic_vector(4 downto 0);
        ADC2_MODE       : in     vl_logic_vector(3 downto 0);
        ADC2_TVC        : in     vl_logic_vector(7 downto 0);
        ADC2_STC        : in     vl_logic_vector(7 downto 0);
        ADC2_ADCSTART   : in     vl_logic;
        ACB_RST         : in     vl_logic;
        ACB_WEN         : in     vl_logic;
        ACB_ADDR        : in     vl_logic_vector(7 downto 0);
        ACB_WDATA       : in     vl_logic_vector(7 downto 0);
        ADC_VAREFOUT    : out    vl_logic;
        ACB_RDATA       : out    vl_logic_vector(7 downto 0);
        ADC0_BUSY       : out    vl_logic;
        ADC0_CALIBRATE  : out    vl_logic;
        ADC0_DATAVALID  : out    vl_logic;
        ADC0_SAMPLE     : out    vl_logic;
        ADC0_RESULT     : out    vl_logic_vector(11 downto 0);
        ADC1_BUSY       : out    vl_logic;
        ADC1_CALIBRATE  : out    vl_logic;
        ADC1_DATAVALID  : out    vl_logic;
        ADC1_SAMPLE     : out    vl_logic;
        ADC1_RESULT     : out    vl_logic_vector(11 downto 0);
        ADC2_BUSY       : out    vl_logic;
        ADC2_CALIBRATE  : out    vl_logic;
        ADC2_DATAVALID  : out    vl_logic;
        ADC2_SAMPLE     : out    vl_logic;
        ADC2_RESULT     : out    vl_logic_vector(11 downto 0);
        DACOUT0         : out    vl_logic;
        DACOUT1         : out    vl_logic;
        DACOUT2         : out    vl_logic;
        DIG_ADC         : out    vl_logic_vector(11 downto 0);
        OBD_DIN         : in     vl_logic_vector(2 downto 0);
        OBD_CLKIN       : in     vl_logic_vector(2 downto 0);
        OBD_ENABLE      : in     vl_logic_vector(2 downto 0);
        COMPARATOR      : out    vl_logic_vector(11 downto 0)
    );
end F2AB;
