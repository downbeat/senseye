// ********************************************************************/
// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//
// Description:	CoreAHBLite - user testbench
//
// Revision Information:
// Date			Description
// ----			-----------------------------------------
// 10Feb10		Production Release Version 3.1
//
// SVN Revision Information:
// SVN $Revision: 3935 $
// SVN $Date: 2008-10-30 18:43:44 -0700 (Thu, 30 Oct 2008) $
//
// Resolved SARs
// SAR      Date     Who   Description
//
// Notes:
// 1. best viewed with tabstops set to "4" (tabs used throughout file)
//
// *********************************************************************/

`timescale 1ns/1ps

module testbench();

// location of this can be overridden at compile time (+incdir switch)
//`include "../../../../coreparameters.v"
`include "coreparameters.v"

parameter SYSCLK_PERIOD = 10; // 100MHz

// the locations and names of these can be overridden at run time
parameter MASTER0_VECTFILE	= "coreahblite_usertb_ahb_master0.vec";
parameter MASTER1_VECTFILE	= "coreahblite_usertb_ahb_master1.vec";

// propagation delay in ns
parameter TPD			= 3;

reg					stopsim=0;
  
reg					SYSCLK;
reg					SYSRSTN;
// using HCLK & HRESETN from master 0 to connect to CoreAHBLite
wire				HCLK;
wire				HRESETN;

// control remap signal from master 0 BFM
wire				REMAP_M0;

// GPIO for 2 master BFM's
wire	[31:0]		GP_OUT_M0;
wire	[31:0]		GP_OUT_M1;
// GP_IN shared
wire	[31:0]		GP_IN;

// signals for testbench request/acknowledgement between masters
wire				M0_REQ;
wire				M0_ACK;
wire				M1_REQ;
wire				M1_ACK;


wire				HREADY_M0;
wire	[1:0]		HRESP_M0;
wire	[31:0]		HRDATA_M0;
wire	[1:0]		HTRANS_M0;
wire	[2:0]		HSIZE_M0;
wire				HWRITE_M0;
wire				HMASTLOCK_M0;
wire	[31:0]		HADDR_M0;
wire	[31:0]		HWDATA_M0;
wire	[2:0]		HBURST_M0;
wire	[3:0]		HPROT_M0;

wire				HREADY_M1;
wire	[1:0]		HRESP_M1;
wire	[31:0]		HRDATA_M1;
wire	[1:0]		HTRANS_M1;
wire	[2:0]		HSIZE_M1;
wire				HWRITE_M1;
wire				HMASTLOCK_M1;
wire	[31:0]		HADDR_M1;
wire	[31:0]		HWDATA_M1;
wire	[2:0]		HBURST_M1;
wire	[3:0]		HPROT_M1;

wire				HWRITE_S0;
wire	[2:0]		HSIZE_S0;
wire	[1:0]		HTRANS_S0;
wire	[31:0]		HWDATA_S0;
wire				HREADYIN_S0;
wire				HSEL_S0;
wire	[31:0]		HADDR_S0;
wire	[31:0]		HRDATA_S0;
wire	[1:0]		HRESP_S0;
wire				HREADY_S0;
wire				HMASTLOCK_S0;
wire	[2:0]		HBURST_S0;
wire	[3:0]		HPROT_S0;

wire				HWRITE_S1;
wire	[2:0]		HSIZE_S1;
wire	[1:0]		HTRANS_S1;
wire	[31:0]		HWDATA_S1;
wire				HREADYIN_S1;
wire				HSEL_S1;
wire	[31:0]		HADDR_S1;
wire	[31:0]		HRDATA_S1;
wire	[1:0]		HRESP_S1;
wire				HREADY_S1;
wire				HMASTLOCK_S1;
wire	[2:0]		HBURST_S1;
wire	[3:0]		HPROT_S1;

wire				HWRITE_S2;
wire	[2:0]		HSIZE_S2;
wire	[1:0]		HTRANS_S2;
wire	[31:0]		HWDATA_S2;
wire				HREADYIN_S2;
wire				HSEL_S2;
wire	[31:0]		HADDR_S2;
wire	[31:0]		HRDATA_S2;
wire	[1:0]		HRESP_S2;
wire				HREADY_S2;
wire				HMASTLOCK_S2;
wire	[2:0]		HBURST_S2;
wire	[3:0]		HPROT_S2;

wire				HWRITE_S3;
wire	[2:0]		HSIZE_S3;
wire	[1:0]		HTRANS_S3;
wire	[31:0]		HWDATA_S3;
wire				HREADYIN_S3;
wire				HSEL_S3;
wire	[31:0]		HADDR_S3;
wire	[31:0]		HRDATA_S3;
wire	[1:0]		HRESP_S3;
wire				HREADY_S3;
wire				HMASTLOCK_S3;
wire	[2:0]		HBURST_S3;
wire	[3:0]		HPROT_S3;

wire				HWRITE_S4;
wire	[2:0]		HSIZE_S4;
wire	[1:0]		HTRANS_S4;
wire	[31:0]		HWDATA_S4;
wire				HREADYIN_S4;
wire				HSEL_S4;
wire	[31:0]		HADDR_S4;
wire	[31:0]		HRDATA_S4;
wire	[1:0]		HRESP_S4;
wire				HREADY_S4;
wire				HMASTLOCK_S4;
wire	[2:0]		HBURST_S4;
wire	[3:0]		HPROT_S4;

wire				HWRITE_S5;
wire	[2:0]		HSIZE_S5;
wire	[1:0]		HTRANS_S5;
wire	[31:0]		HWDATA_S5;
wire				HREADYIN_S5;
wire				HSEL_S5;
wire	[31:0]		HADDR_S5;
wire	[31:0]		HRDATA_S5;
wire	[1:0]		HRESP_S5;
wire				HREADY_S5;
wire				HMASTLOCK_S5;
wire	[2:0]		HBURST_S5;
wire	[3:0]		HPROT_S5;

wire				HWRITE_S6;
wire	[2:0]		HSIZE_S6;
wire	[1:0]		HTRANS_S6;
wire	[31:0]		HWDATA_S6;
wire				HREADYIN_S6;
wire				HSEL_S6;
wire	[31:0]		HADDR_S6;
wire	[31:0]		HRDATA_S6;
wire	[1:0]		HRESP_S6;
wire				HREADY_S6;
wire				HMASTLOCK_S6;
wire	[2:0]		HBURST_S6;
wire	[3:0]		HPROT_S6;

wire				HWRITE_S7;
wire	[2:0]		HSIZE_S7;
wire	[1:0]		HTRANS_S7;
wire	[31:0]		HWDATA_S7;
wire				HREADYIN_S7;
wire				HSEL_S7;
wire	[31:0]		HADDR_S7;
wire	[31:0]		HRDATA_S7;
wire	[1:0]		HRESP_S7;
wire				HREADY_S7;
wire				HMASTLOCK_S7;
wire	[2:0]		HBURST_S7;
wire	[3:0]		HPROT_S7;

wire				HWRITE_S8;
wire	[2:0]		HSIZE_S8;
wire	[1:0]		HTRANS_S8;
wire	[31:0]		HWDATA_S8;
wire				HREADYIN_S8;
wire				HSEL_S8;
wire	[31:0]		HADDR_S8;
wire	[31:0]		HRDATA_S8;
wire	[1:0]		HRESP_S8;
wire				HREADY_S8;
wire				HMASTLOCK_S8;
wire	[2:0]		HBURST_S8;
wire	[3:0]		HPROT_S8;

wire				HWRITE_S9;
wire	[2:0]		HSIZE_S9;
wire	[1:0]		HTRANS_S9;
wire	[31:0]		HWDATA_S9;
wire				HREADYIN_S9;
wire				HSEL_S9;
wire	[31:0]		HADDR_S9;
wire	[31:0]		HRDATA_S9;
wire	[1:0]		HRESP_S9;
wire				HREADY_S9;
wire				HMASTLOCK_S9;
wire	[2:0]		HBURST_S9;
wire	[3:0]		HPROT_S9;

wire				HWRITE_S10;
wire	[2:0]		HSIZE_S10;
wire	[1:0]		HTRANS_S10;
wire	[31:0]		HWDATA_S10;
wire				HREADYIN_S10;
wire				HSEL_S10;
wire	[31:0]		HADDR_S10;
wire	[31:0]		HRDATA_S10;
wire	[1:0]		HRESP_S10;
wire				HREADY_S10;
wire				HMASTLOCK_S10;
wire	[2:0]		HBURST_S10;
wire	[3:0]		HPROT_S10;

wire				HWRITE_S11;
wire	[2:0]		HSIZE_S11;
wire	[1:0]		HTRANS_S11;
wire	[31:0]		HWDATA_S11;
wire				HREADYIN_S11;
wire				HSEL_S11;
wire	[31:0]		HADDR_S11;
wire	[31:0]		HRDATA_S11;
wire	[1:0]		HRESP_S11;
wire				HREADY_S11;
wire				HMASTLOCK_S11;
wire	[2:0]		HBURST_S11;
wire	[3:0]		HPROT_S11;

wire				HWRITE_S12;
wire	[2:0]		HSIZE_S12;
wire	[1:0]		HTRANS_S12;
wire	[31:0]		HWDATA_S12;
wire				HREADYIN_S12;
wire				HSEL_S12;
wire	[31:0]		HADDR_S12;
wire	[31:0]		HRDATA_S12;
wire	[1:0]		HRESP_S12;
wire				HREADY_S12;
wire				HMASTLOCK_S12;
wire	[2:0]		HBURST_S12;
wire	[3:0]		HPROT_S12;

wire				HWRITE_S13;
wire	[2:0]		HSIZE_S13;
wire	[1:0]		HTRANS_S13;
wire	[31:0]		HWDATA_S13;
wire				HREADYIN_S13;
wire				HSEL_S13;
wire	[31:0]		HADDR_S13;
wire	[31:0]		HRDATA_S13;
wire	[1:0]		HRESP_S13;
wire				HREADY_S13;
wire				HMASTLOCK_S13;
wire	[2:0]		HBURST_S13;
wire	[3:0]		HPROT_S13;

wire				HWRITE_S14;
wire	[2:0]		HSIZE_S14;
wire	[1:0]		HTRANS_S14;
wire	[31:0]		HWDATA_S14;
wire				HREADYIN_S14;
wire				HSEL_S14;
wire	[31:0]		HADDR_S14;
wire	[31:0]		HRDATA_S14;
wire	[1:0]		HRESP_S14;
wire				HREADY_S14;
wire				HMASTLOCK_S14;
wire	[2:0]		HBURST_S14;
wire	[3:0]		HPROT_S14;

wire				HWRITE_S15;
wire	[2:0]		HSIZE_S15;
wire	[1:0]		HTRANS_S15;
wire	[31:0]		HWDATA_S15;
wire				HREADYIN_S15;
wire				HSEL_S15;
wire	[31:0]		HADDR_S15;
wire	[31:0]		HRDATA_S15;
wire	[1:0]		HRESP_S15;
wire				HREADY_S15;
wire				HMASTLOCK_S15;
wire	[2:0]		HBURST_S15;
wire	[3:0]		HPROT_S15;

wire				HWRITE_SHG;
wire	[2:0]		HSIZE_SHG;
wire	[1:0]		HTRANS_SHG;
wire	[31:0]		HWDATA_SHG;
wire				HREADYIN_SHG;
wire				HSEL_SHG;
wire	[31:0]		HADDR_SHG;
wire	[31:0]		HRDATA_SHG;
wire	[1:0]		HRESP_SHG;
wire				HREADY_SHG;
wire				HMASTLOCK_SHG;
wire	[2:0]		HBURST_SHG;
wire	[3:0]		HPROT_SHG;

// Init/Config client 0 Signals
wire				INITDATVAL_C0;
wire				INITDONE_C0;
wire	[11:0]		INITADDR_C0;
wire	[31:0]		INITDATA_C0;

// Init/Config client 1 Signals
wire				INITDATVAL_C1;
wire				INITDONE_C1;
wire	[11:0]		INITADDR_C1;
wire	[31:0]		INITDATA_C1;

// Init/Config client 2 Signals
wire				INITDATVAL_C2;
wire				INITDONE_C2;
wire	[11:0]		INITADDR_C2;
wire	[31:0]		INITDATA_C2;

// Init/Config client 3 Signals
wire				INITDATVAL_C3;
wire				INITDONE_C3;
wire	[11:0]		INITADDR_C3;
wire	[31:0]		INITDATA_C3;

// Init/Config client 4 Signals
wire				INITDATVAL_C4;
wire				INITDONE_C4;
wire	[11:0]		INITADDR_C4;
wire	[31:0]		INITDATA_C4;

// Init/Config client 5 Signals
wire				INITDATVAL_C5;
wire				INITDONE_C5;
wire	[11:0]		INITADDR_C5;
wire	[31:0]		INITDATA_C5;

// Init/Config client 6 Signals
wire				INITDATVAL_C6;
wire				INITDONE_C6;
wire	[11:0]		INITADDR_C6;
wire	[31:0]		INITDATA_C6;

// Init/Config client 7 Signals
wire				INITDATVAL_C7;
wire				INITDONE_C7;
wire	[11:0]		INITADDR_C7;
wire	[31:0]		INITDATA_C7;

// Init/Config client 8 Signals
wire				INITDATVAL_C8;
wire				INITDONE_C8;
wire	[11:0]		INITADDR_C8;
wire	[31:0]		INITDATA_C8;

// Init/Config client 9 Signals
wire				INITDATVAL_C9;
wire				INITDONE_C9;
wire	[11:0]		INITADDR_C9;
wire	[31:0]		INITDATA_C9;

// Init/Config client 10 Signals
wire				INITDATVAL_C10;
wire				INITDONE_C10;
wire	[11:0]		INITADDR_C10;
wire	[31:0]		INITDATA_C10;

// Init/Config client 11 Signals
wire				INITDATVAL_C11;
wire				INITDONE_C11;
wire	[11:0]		INITADDR_C11;
wire	[31:0]		INITDATA_C11;

// Init/Config client 12 Signals
wire				INITDATVAL_C12;
wire				INITDONE_C12;
wire	[11:0]		INITADDR_C12;
wire	[31:0]		INITDATA_C12;

// Init/Config client 13 Signals
wire				INITDATVAL_C13;
wire				INITDONE_C13;
wire	[11:0]		INITADDR_C13;
wire	[31:0]		INITDATA_C13;

// Init/Config client 14 Signals
wire				INITDATVAL_C14;
wire				INITDONE_C14;
wire	[11:0]		INITADDR_C14;
wire	[31:0]		INITDATA_C14;

// Init/Config client 15 Signals
wire				INITDATVAL_C15;
wire				INITDONE_C15;
wire	[11:0]		INITADDR_C15;
wire	[31:0]		INITDATA_C15;





wire				FINISHED_master0;
wire				FINISHED_master1;

initial
begin
    SYSCLK = 1'b0;
    SYSRSTN = 1'b0;

	// Release system reset
    #(SYSCLK_PERIOD * 4)
        SYSRSTN = 1'b1;

	// wait until both BFM's are finished
	while (!((FINISHED_master0===1'b1) && (FINISHED_master1===1'b1)))
	begin
		@ (posedge SYSCLK); #TPD;
	end
	stopsim=1;
	#1;
	$stop;
end

// tie-off unused inputs to DUT
assign HBURST_M0	= 3'b0;
assign HBURST_M1	= 3'b0;
assign HPROT_M0		= 4'b0;
assign HPROT_M1		= 4'b0;
assign HRESP_S0[1]	= 1'b0;
assign HRESP_S1[1]	= 1'b0;
assign HRESP_S2[1]	= 1'b0;
assign HRESP_S3[1]	= 1'b0;
assign HRESP_S4[1]	= 1'b0;
assign HRESP_S5[1]	= 1'b0;
assign HRESP_S6[1]	= 1'b0;
assign HRESP_S7[1]	= 1'b0;
assign HRESP_S8[1]	= 1'b0;
assign HRESP_S9[1]	= 1'b0;
assign HRESP_S10[1]	= 1'b0;
assign HRESP_S11[1]	= 1'b0;
assign HRESP_S12[1]	= 1'b0;
assign HRESP_S13[1]	= 1'b0;
assign HRESP_S14[1]	= 1'b0;
assign HRESP_S15[1]	= 1'b0;
assign HRESP_SHG[1]	= 1'b0;

// SYSCLK signal
always @(SYSCLK)
    #(SYSCLK_PERIOD / 2)
    SYSCLK <= !SYSCLK;

// Instantiate module to test
CoreAHBLite #( 
	.FAMILY(FAMILY),
	.MODE_CFG(MODE_CFG),
	.M0_AHBSLOT0ENABLE(M0_AHBSLOT0ENABLE),
	.M0_AHBSLOT1ENABLE(M0_AHBSLOT1ENABLE ),
	.M0_AHBSLOT2ENABLE(M0_AHBSLOT2ENABLE ),
	.M0_AHBSLOT3ENABLE(M0_AHBSLOT3ENABLE ),
	.M0_AHBSLOT4ENABLE(M0_AHBSLOT4ENABLE ),
	.M0_AHBSLOT5ENABLE(M0_AHBSLOT5ENABLE ),
	.M0_AHBSLOT6ENABLE(M0_AHBSLOT6ENABLE ),
	.M0_AHBSLOT7ENABLE(M0_AHBSLOT7ENABLE ),
	.M0_AHBSLOT8ENABLE(M0_AHBSLOT8ENABLE ),
	.M0_AHBSLOT9ENABLE(M0_AHBSLOT9ENABLE ),
	.M0_AHBSLOT10ENABLE(M0_AHBSLOT10ENABLE),
	.M0_AHBSLOT11ENABLE(M0_AHBSLOT11ENABLE),
	.M0_AHBSLOT12ENABLE(M0_AHBSLOT12ENABLE),
	.M0_AHBSLOT13ENABLE(M0_AHBSLOT13ENABLE),
	.M0_AHBSLOT14ENABLE(M0_AHBSLOT14ENABLE),
	.M0_AHBSLOT15ENABLE(M0_AHBSLOT15ENABLE),
	.M1_AHBSLOT0ENABLE(M1_AHBSLOT0ENABLE ),
	.M1_AHBSLOT1ENABLE(M1_AHBSLOT1ENABLE ),
	.M1_AHBSLOT2ENABLE(M1_AHBSLOT2ENABLE ),
	.M1_AHBSLOT3ENABLE(M1_AHBSLOT3ENABLE ),
	.M1_AHBSLOT4ENABLE(M1_AHBSLOT4ENABLE ),
	.M1_AHBSLOT5ENABLE(M1_AHBSLOT5ENABLE ),
	.M1_AHBSLOT6ENABLE(M1_AHBSLOT6ENABLE ),
	.M1_AHBSLOT7ENABLE(M1_AHBSLOT7ENABLE ),
	.M1_AHBSLOT8ENABLE(M1_AHBSLOT8ENABLE ),
	.M1_AHBSLOT9ENABLE(M1_AHBSLOT9ENABLE ),
	.M1_AHBSLOT10ENABLE(M1_AHBSLOT10ENABLE),
	.M1_AHBSLOT11ENABLE(M1_AHBSLOT11ENABLE),
	.M1_AHBSLOT12ENABLE(M1_AHBSLOT12ENABLE),
	.M1_AHBSLOT13ENABLE(M1_AHBSLOT13ENABLE),
	.M1_AHBSLOT14ENABLE(M1_AHBSLOT14ENABLE),
	.M1_AHBSLOT15ENABLE(M1_AHBSLOT15ENABLE),
	.M0_HUGESLOTENABLE(M0_HUGESLOTENABLE),
	.M1_HUGESLOTENABLE(M1_HUGESLOTENABLE),
	.HADDR_SHG_CFG(HADDR_SHG_CFG),
	.M0_INITCFG0ENABLE(M0_INITCFG0ENABLE),
	.M0_INITCFG1ENABLE(M0_INITCFG1ENABLE),
	.M0_INITCFG2ENABLE(M0_INITCFG2ENABLE),
	.M0_INITCFG3ENABLE(M0_INITCFG3ENABLE),
	.M0_INITCFG4ENABLE(M0_INITCFG4ENABLE),
	.M0_INITCFG5ENABLE(M0_INITCFG5ENABLE),
	.M0_INITCFG6ENABLE(M0_INITCFG6ENABLE),
	.M0_INITCFG7ENABLE(M0_INITCFG7ENABLE),
	.M0_INITCFG8ENABLE(M0_INITCFG8ENABLE),
	.M0_INITCFG9ENABLE(M0_INITCFG9ENABLE),
	.M0_INITCFG10ENABLE(M0_INITCFG10ENABLE),
	.M0_INITCFG11ENABLE(M0_INITCFG11ENABLE),
	.M0_INITCFG12ENABLE(M0_INITCFG12ENABLE),
	.M0_INITCFG13ENABLE(M0_INITCFG13ENABLE),
	.M0_INITCFG14ENABLE(M0_INITCFG14ENABLE),
	.M0_INITCFG15ENABLE(M0_INITCFG15ENABLE),
	.M1_INITCFG0ENABLE(M1_INITCFG0ENABLE),
	.M1_INITCFG1ENABLE(M1_INITCFG1ENABLE),
	.M1_INITCFG2ENABLE(M1_INITCFG2ENABLE),
	.M1_INITCFG3ENABLE(M1_INITCFG3ENABLE),
	.M1_INITCFG4ENABLE(M1_INITCFG4ENABLE),
	.M1_INITCFG5ENABLE(M1_INITCFG5ENABLE),
	.M1_INITCFG6ENABLE(M1_INITCFG6ENABLE),
	.M1_INITCFG7ENABLE(M1_INITCFG7ENABLE),
	.M1_INITCFG8ENABLE(M1_INITCFG8ENABLE),
	.M1_INITCFG9ENABLE(M1_INITCFG9ENABLE),
	.M1_INITCFG10ENABLE(M1_INITCFG10ENABLE),
	.M1_INITCFG11ENABLE(M1_INITCFG11ENABLE),
	.M1_INITCFG12ENABLE(M1_INITCFG12ENABLE),
	.M1_INITCFG13ENABLE(M1_INITCFG13ENABLE),
	.M1_INITCFG14ENABLE(M1_INITCFG14ENABLE),
	.M1_INITCFG15ENABLE(M1_INITCFG15ENABLE)
) u_coreahblite (
	// ResetController interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),

	// controls master 0 memory aliasing (swaps slots 0 and 1)
	.REMAP_M0(REMAP_M0),

	// Mirrored master AHB-Lite interface to Master 0
	// Inputs
	.HADDR_M0(HADDR_M0),
	.HMASTLOCK_M0(HMASTLOCK_M0),
	.HSIZE_M0(HSIZE_M0),
	.HTRANS_M0(HTRANS_M0),
	.HWRITE_M0(HWRITE_M0),
	.HWDATA_M0(HWDATA_M0),
	.HBURST_M0(HBURST_M0),
	.HPROT_M0(HPROT_M0),
	// Outputs
	.HRESP_M0(HRESP_M0),
	.HRDATA_M0(HRDATA_M0),
	.HREADY_M0(HREADY_M0),

	// Mirrored master AHB-Lite interface to Master 1
	// Inputs
	.HADDR_M1(HADDR_M1),
	.HMASTLOCK_M1(HMASTLOCK_M1),
	.HSIZE_M1(HSIZE_M1),
	.HTRANS_M1(HTRANS_M1),
	.HWRITE_M1(HWRITE_M1),
	.HWDATA_M1(HWDATA_M1),
	.HBURST_M1(HBURST_M1),
	.HPROT_M1(HPROT_M1),

	// Outputs
	.HRESP_M1(HRESP_M1),
	.HRDATA_M1(HRDATA_M1),
	.HREADY_M1(HREADY_M1),

	// Mirrored slave AHB-Lite interface to Slave 0
	// Inputs
	.HRDATA_S0(HRDATA_S0),
	.HREADYOUT_S0(HREADY_S0),
	.HRESP_S0(HRESP_S0),
	// Outputs
	.HSEL_S0(HSEL_S0),
	.HADDR_S0(HADDR_S0),
	.HSIZE_S0(HSIZE_S0),
	.HTRANS_S0(HTRANS_S0),
	.HWRITE_S0(HWRITE_S0),
	.HWDATA_S0(HWDATA_S0),
	.HREADY_S0(HREADYIN_S0),
	.HMASTLOCK_S0(HMASTLOCK_S0),
	.HBURST_S0(HBURST_S0),
	.HPROT_S0(HPROT_S0),

	// Mirrored slave AHB-Lite interface to Slave 1
	// Inputs
	.HRDATA_S1(HRDATA_S1),
	.HREADYOUT_S1(HREADY_S1),
	.HRESP_S1(HRESP_S1),
	// Outputs
	.HSEL_S1(HSEL_S1),
	.HADDR_S1(HADDR_S1),
	.HSIZE_S1(HSIZE_S1),
	.HTRANS_S1(HTRANS_S1),
	.HWRITE_S1(HWRITE_S1),
	.HWDATA_S1(HWDATA_S1),
	.HREADY_S1(HREADYIN_S1),
	.HMASTLOCK_S1(HMASTLOCK_S1),
	.HBURST_S1(HBURST_S1),
	.HPROT_S1(HPROT_S1),

	// Mirrored slave AHB-Lite interface to Slave 2
	// Inputs
	.HRDATA_S2(HRDATA_S2),
	.HREADYOUT_S2(HREADY_S2),
	.HRESP_S2(HRESP_S2),
	// Outputs
	.HSEL_S2(HSEL_S2),
	.HADDR_S2(HADDR_S2),
	.HSIZE_S2(HSIZE_S2),
	.HTRANS_S2(HTRANS_S2),
	.HWRITE_S2(HWRITE_S2),
	.HWDATA_S2(HWDATA_S2),
	.HREADY_S2(HREADYIN_S2),
	.HMASTLOCK_S2(HMASTLOCK_S2),
	.HBURST_S2(HBURST_S2),
	.HPROT_S2(HPROT_S2),

	// Mirrored slave AHB-Lite interface to Slave 3
	// Inputs
	.HRDATA_S3(HRDATA_S3),
	.HREADYOUT_S3(HREADY_S3),
	.HRESP_S3(HRESP_S3),
	// Output
	.HSEL_S3(HSEL_S3),
	.HADDR_S3(HADDR_S3),
	.HSIZE_S3(HSIZE_S3),
	.HTRANS_S3(HTRANS_S3),
	.HWRITE_S3(HWRITE_S3),
	.HWDATA_S3(HWDATA_S3),
	.HREADY_S3(HREADYIN_S3),
	.HMASTLOCK_S3(HMASTLOCK_S3),
	.HBURST_S3(HBURST_S3),
	.HPROT_S3(HPROT_S3),

	// Mirrored slave AHB-Lite interface to Slave 4
	// Inputs
	.HRDATA_S4(HRDATA_S4),
	.HREADYOUT_S4(HREADY_S4),
	.HRESP_S4(HRESP_S4),
	// Output
	.HSEL_S4(HSEL_S4),
	.HADDR_S4(HADDR_S4),
	.HSIZE_S4(HSIZE_S4),
	.HTRANS_S4(HTRANS_S4),
	.HWRITE_S4(HWRITE_S4),
	.HWDATA_S4(HWDATA_S4),
	.HREADY_S4(HREADYIN_S4),
	.HMASTLOCK_S4(HMASTLOCK_S4),
	.HBURST_S4(HBURST_S4),
	.HPROT_S4(HPROT_S4),

	// Mirrored slave AHB-Lite interface to Slave 5
	// Inputs
	.HRDATA_S5(HRDATA_S5),
	.HREADYOUT_S5(HREADY_S5),
	.HRESP_S5(HRESP_S5),
	// Output
	.HSEL_S5(HSEL_S5),
	.HADDR_S5(HADDR_S5),
	.HSIZE_S5(HSIZE_S5),
	.HTRANS_S5(HTRANS_S5),
	.HWRITE_S5(HWRITE_S5),
	.HWDATA_S5(HWDATA_S5),
	.HREADY_S5(HREADYIN_S5),
	.HMASTLOCK_S5(HMASTLOCK_S5),
	.HBURST_S5(HBURST_S5),
	.HPROT_S5(HPROT_S5),

	// Mirrored slave AHB-Lite interface to Slave 6
	// Inputs
	.HRDATA_S6(HRDATA_S6),
	.HREADYOUT_S6(HREADY_S6),
	.HRESP_S6(HRESP_S6),
	// Output
	.HSEL_S6(HSEL_S6),
	.HADDR_S6(HADDR_S6),
	.HSIZE_S6(HSIZE_S6),
	.HTRANS_S6(HTRANS_S6),
	.HWRITE_S6(HWRITE_S6),
	.HWDATA_S6(HWDATA_S6),
	.HREADY_S6(HREADYIN_S6),
	.HMASTLOCK_S6(HMASTLOCK_S6),
	.HBURST_S6(HBURST_S6),
	.HPROT_S6(HPROT_S6),

	// Mirrored slave AHB-Lite interface to Slave 7
	// Inputs
	.HRDATA_S7(HRDATA_S7),
	.HREADYOUT_S7(HREADY_S7),
	.HRESP_S7(HRESP_S7),
	// Output
	.HSEL_S7(HSEL_S7),
	.HADDR_S7(HADDR_S7),
	.HSIZE_S7(HSIZE_S7),
	.HTRANS_S7(HTRANS_S7),
	.HWRITE_S7(HWRITE_S7),
	.HWDATA_S7(HWDATA_S7),
	.HREADY_S7(HREADYIN_S7),
	.HMASTLOCK_S7(HMASTLOCK_S7),
	.HBURST_S7(HBURST_S7),
	.HPROT_S7(HPROT_S7),

	// Mirrored slave AHB-Lite interface to Slave 8
	// Inputs
	.HRDATA_S8(HRDATA_S8),
	.HREADYOUT_S8(HREADY_S8),
	.HRESP_S8(HRESP_S8),
	// Output
	.HSEL_S8(HSEL_S8),
	.HADDR_S8(HADDR_S8),
	.HSIZE_S8(HSIZE_S8),
	.HTRANS_S8(HTRANS_S8),
	.HWRITE_S8(HWRITE_S8),
	.HWDATA_S8(HWDATA_S8),
	.HREADY_S8(HREADYIN_S8),
	.HMASTLOCK_S8(HMASTLOCK_S8),
	.HBURST_S8(HBURST_S8),
	.HPROT_S8(HPROT_S8),

	// Mirrored slave AHB-Lite interface to Slave 9
	// Inputs
	.HRDATA_S9(HRDATA_S9),
	.HREADYOUT_S9(HREADY_S9),
	.HRESP_S9(HRESP_S9),
	// Output
	.HSEL_S9(HSEL_S9),
	.HADDR_S9(HADDR_S9),
	.HSIZE_S9(HSIZE_S9),
	.HTRANS_S9(HTRANS_S9),
	.HWRITE_S9(HWRITE_S9),
	.HWDATA_S9(HWDATA_S9),
	.HREADY_S9(HREADYIN_S9),
	.HMASTLOCK_S9(HMASTLOCK_S9),
	.HBURST_S9(HBURST_S9),
	.HPROT_S9(HPROT_S9),

	// Mirrored slave AHB-Lite interface to Slave 10
	// Inputs
	.HRDATA_S10(HRDATA_S10),
	.HREADYOUT_S10(HREADY_S10),
	.HRESP_S10(HRESP_S10),
	// Output
	.HSEL_S10(HSEL_S10),
	.HADDR_S10(HADDR_S10),
	.HSIZE_S10(HSIZE_S10),
	.HTRANS_S10(HTRANS_S10),
	.HWRITE_S10(HWRITE_S10),
	.HWDATA_S10(HWDATA_S10),
	.HREADY_S10(HREADYIN_S10),
	.HMASTLOCK_S10(HMASTLOCK_S10),
	.HBURST_S10(HBURST_S10),
	.HPROT_S10(HPROT_S10),

	// Mirrored slave AHB-Lite interface to Slave 11
	// Inputs
	.HRDATA_S11(HRDATA_S11),
	.HREADYOUT_S11(HREADY_S11),
	.HRESP_S11(HRESP_S11),
	// Output
	.HSEL_S11(HSEL_S11),
	.HADDR_S11(HADDR_S11),
	.HSIZE_S11(HSIZE_S11),
	.HTRANS_S11(HTRANS_S11),
	.HWRITE_S11(HWRITE_S11),
	.HWDATA_S11(HWDATA_S11),
	.HREADY_S11(HREADYIN_S11),
	.HMASTLOCK_S11(HMASTLOCK_S11),
	.HBURST_S11(HBURST_S11),
	.HPROT_S11(HPROT_S11),

	// Mirrored slave AHB-Lite interface to Slave 12
	// Inputs
	.HRDATA_S12(HRDATA_S12),
	.HREADYOUT_S12(HREADY_S12),
	.HRESP_S12(HRESP_S12),
	// Output
	.HSEL_S12(HSEL_S12),
	.HADDR_S12(HADDR_S12),
	.HSIZE_S12(HSIZE_S12),
	.HTRANS_S12(HTRANS_S12),
	.HWRITE_S12(HWRITE_S12),
	.HWDATA_S12(HWDATA_S12),
	.HREADY_S12(HREADYIN_S12),
	.HMASTLOCK_S12(HMASTLOCK_S12),
	.HBURST_S12(HBURST_S12),
	.HPROT_S12(HPROT_S12),

	// Mirrored slave AHB-Lite interface to Slave 13
	// Inputs
	.HRDATA_S13(HRDATA_S13),
	.HREADYOUT_S13(HREADY_S13),
	.HRESP_S13(HRESP_S13),
	// Output
	.HSEL_S13(HSEL_S13),
	.HADDR_S13(HADDR_S13),
	.HSIZE_S13(HSIZE_S13),
	.HTRANS_S13(HTRANS_S13),
	.HWRITE_S13(HWRITE_S13),
	.HWDATA_S13(HWDATA_S13),
	.HREADY_S13(HREADYIN_S13),
	.HMASTLOCK_S13(HMASTLOCK_S13),
	.HBURST_S13(HBURST_S13),
	.HPROT_S13(HPROT_S13),

	// Mirrored slave AHB-Lite interface to Slave 14
	// Inputs
	.HRDATA_S14(HRDATA_S14),
	.HREADYOUT_S14(HREADY_S14),
	.HRESP_S14(HRESP_S14),
	// Output
	.HSEL_S14(HSEL_S14),
	.HADDR_S14(HADDR_S14),
	.HSIZE_S14(HSIZE_S14),
	.HTRANS_S14(HTRANS_S14),
	.HWRITE_S14(HWRITE_S14),
	.HWDATA_S14(HWDATA_S14),
	.HREADY_S14(HREADYIN_S14),
	.HMASTLOCK_S14(HMASTLOCK_S14),
	.HBURST_S14(HBURST_S14),
	.HPROT_S14(HPROT_S14),

	// Mirrored slave AHB-Lite interface to Slave 15
	// Inputs
	.HRDATA_S15(HRDATA_S15),
	.HREADYOUT_S15(HREADY_S15),
	.HRESP_S15(HRESP_S15),
	// Output
	.HSEL_S15(HSEL_S15),
	.HADDR_S15(HADDR_S15),
	.HSIZE_S15(HSIZE_S15),
	.HTRANS_S15(HTRANS_S15),
	.HWRITE_S15(HWRITE_S15),
	.HWDATA_S15(HWDATA_S15),
	.HREADY_S15(HREADYIN_S15),
	.HMASTLOCK_S15(HMASTLOCK_S15),
	.HBURST_S15(HBURST_S15),
	.HPROT_S15(HPROT_S15),

	// Mirrored slave AHB-Lite interface to Huge Slave
	// Inputs
	.HRDATA_SHG(HRDATA_SHG),
	.HREADYOUT_SHG(HREADY_SHG),
	.HRESP_SHG(HRESP_SHG),
	// Outputs
	.HSEL_SHG(HSEL_SHG),
	.HADDR_SHG(HADDR_SHG),
	.HSIZE_SHG(HSIZE_SHG),
	.HTRANS_SHG(HTRANS_SHG),
	.HWRITE_SHG(HWRITE_SHG),
	.HWDATA_SHG(HWDATA_SHG),
	.HREADY_SHG(HREADYIN_SHG),
	.HMASTLOCK_SHG(HMASTLOCK_SHG),
	.HBURST_SHG(HBURST_SHG),
	.HPROT_SHG(HPROT_SHG),

	// outputs to Init/Config clients
	.INITDATVAL_C0(INITDATVAL_C0),
	.INITDONE_C0(INITDONE_C0),
	.INITADDR_C0(INITADDR_C0),
	.INITDATA_C0(INITDATA_C0),
	.INITDATVAL_C1(INITDATVAL_C1),
	.INITDONE_C1(INITDONE_C1),
	.INITADDR_C1(INITADDR_C1),
	.INITDATA_C1(INITDATA_C1),
	.INITDATVAL_C2(INITDATVAL_C2),
	.INITDONE_C2(INITDONE_C2),
	.INITADDR_C2(INITADDR_C2),
	.INITDATA_C2(INITDATA_C2),
	.INITDATVAL_C3(INITDATVAL_C3),
	.INITDONE_C3(INITDONE_C3),
	.INITADDR_C3(INITADDR_C3),
	.INITDATA_C3(INITDATA_C3),
	.INITDATVAL_C4(INITDATVAL_C4),
	.INITDONE_C4(INITDONE_C4),
	.INITADDR_C4(INITADDR_C4),
	.INITDATA_C4(INITDATA_C4),
	.INITDATVAL_C5(INITDATVAL_C5),
	.INITDONE_C5(INITDONE_C5),
	.INITADDR_C5(INITADDR_C5),
	.INITDATA_C5(INITDATA_C5),
	.INITDATVAL_C6(INITDATVAL_C6),
	.INITDONE_C6(INITDONE_C6),
	.INITADDR_C6(INITADDR_C6),
	.INITDATA_C6(INITDATA_C6),
	.INITDATVAL_C7(INITDATVAL_C7),
	.INITDONE_C7(INITDONE_C7),
	.INITADDR_C7(INITADDR_C7),
	.INITDATA_C7(INITDATA_C7),
	.INITDATVAL_C8(INITDATVAL_C8),
	.INITDONE_C8(INITDONE_C8),
	.INITADDR_C8(INITADDR_C8),
	.INITDATA_C8(INITDATA_C8),
	.INITDATVAL_C9(INITDATVAL_C9),
	.INITDONE_C9(INITDONE_C9),
	.INITADDR_C9(INITADDR_C9),
	.INITDATA_C9(INITDATA_C9),
	.INITDATVAL_C10(INITDATVAL_C10),
	.INITDONE_C10(INITDONE_C10),
	.INITADDR_C10(INITADDR_C10),
	.INITDATA_C10(INITDATA_C10),
	.INITDATVAL_C11(INITDATVAL_C11),
	.INITDONE_C11(INITDONE_C11),
	.INITADDR_C11(INITADDR_C11),
	.INITDATA_C11(INITDATA_C11),
	.INITDATVAL_C12(INITDATVAL_C12),
	.INITDONE_C12(INITDONE_C12),
	.INITADDR_C12(INITADDR_C12),
	.INITDATA_C12(INITDATA_C12),
	.INITDATVAL_C13(INITDATVAL_C13),
	.INITDONE_C13(INITDONE_C13),
	.INITADDR_C13(INITADDR_C13),
	.INITDATA_C13(INITDATA_C13),
	.INITDATVAL_C14(INITDATVAL_C14),
	.INITDONE_C14(INITDONE_C14),
	.INITADDR_C14(INITADDR_C14),
	.INITDATA_C14(INITDATA_C14),
	.INITDATVAL_C15(INITDATVAL_C15),
	.INITDONE_C15(INITDONE_C15),
	.INITADDR_C15(INITADDR_C15),
	.INITDATA_C15(INITDATA_C15)
);

// BFM masters monitor various signals
assign GP_IN = {
	12'b0,
	M1_ACK,
	M1_REQ,
	M0_ACK,
	M0_REQ,
	15'b0,
	REMAP_M0
};


// master 0 BFM
BFM_AHBL #(
	.VECTFILE(MASTER0_VECTFILE),
	// passing testbench parameters to BFM ARGVALUE* parameters
	.ARGVALUE0(FAMILY),
	.ARGVALUE1(MODE_CFG),
	.ARGVALUE2(M0_AHBSLOT0ENABLE),
	.ARGVALUE3(M0_AHBSLOT1ENABLE),
	.ARGVALUE4(M0_AHBSLOT2ENABLE),
	.ARGVALUE5(M0_AHBSLOT3ENABLE),
	.ARGVALUE6(M0_AHBSLOT4ENABLE),
	.ARGVALUE7(M0_AHBSLOT5ENABLE),
	.ARGVALUE8(M0_AHBSLOT6ENABLE),
	.ARGVALUE9(M0_AHBSLOT7ENABLE),
	.ARGVALUE10(M0_AHBSLOT8ENABLE),
	.ARGVALUE11(M0_AHBSLOT9ENABLE),
	.ARGVALUE12(M0_AHBSLOT10ENABLE),
	.ARGVALUE13(M0_AHBSLOT11ENABLE),
	.ARGVALUE14(M0_AHBSLOT12ENABLE),
	.ARGVALUE15(M0_AHBSLOT13ENABLE),
	.ARGVALUE16(M0_AHBSLOT14ENABLE),
	.ARGVALUE17(M0_AHBSLOT15ENABLE),
	.ARGVALUE18(M1_AHBSLOT0ENABLE),
	.ARGVALUE19(M1_AHBSLOT1ENABLE),
	.ARGVALUE20(M1_AHBSLOT2ENABLE),
	.ARGVALUE21(M1_AHBSLOT3ENABLE),
	.ARGVALUE22(M1_AHBSLOT4ENABLE),
	.ARGVALUE23(M1_AHBSLOT5ENABLE),
	.ARGVALUE24(M1_AHBSLOT6ENABLE),
	.ARGVALUE25(M1_AHBSLOT7ENABLE),
	.ARGVALUE26(M1_AHBSLOT8ENABLE),
	.ARGVALUE27(M1_AHBSLOT9ENABLE),
	.ARGVALUE28(M1_AHBSLOT10ENABLE),
	.ARGVALUE29(M1_AHBSLOT11ENABLE),
	.ARGVALUE30(M1_AHBSLOT12ENABLE),
	.ARGVALUE31(M1_AHBSLOT13ENABLE),
	.ARGVALUE32(M1_AHBSLOT14ENABLE),
	.ARGVALUE33(M1_AHBSLOT15ENABLE),
	.ARGVALUE34(M0_HUGESLOTENABLE),
	.ARGVALUE35(M1_HUGESLOTENABLE),
	.ARGVALUE36(HADDR_SHG_CFG),
	.ARGVALUE37(M0_INITCFG0ENABLE),
	.ARGVALUE38(M0_INITCFG1ENABLE),
	.ARGVALUE39(M0_INITCFG2ENABLE),
	.ARGVALUE40(M0_INITCFG3ENABLE),
	.ARGVALUE41(M0_INITCFG4ENABLE),
	.ARGVALUE42(M0_INITCFG5ENABLE),
	.ARGVALUE43(M0_INITCFG6ENABLE),
	.ARGVALUE44(M0_INITCFG7ENABLE),
	.ARGVALUE45(M0_INITCFG8ENABLE),
	.ARGVALUE46(M0_INITCFG9ENABLE),
	.ARGVALUE47(M0_INITCFG10ENABLE),
	.ARGVALUE48(M0_INITCFG11ENABLE),
	.ARGVALUE49(M0_INITCFG12ENABLE),
	.ARGVALUE50(M0_INITCFG13ENABLE),
	.ARGVALUE51(M0_INITCFG14ENABLE),
	.ARGVALUE52(M0_INITCFG15ENABLE),
	.ARGVALUE53(M1_INITCFG0ENABLE),
	.ARGVALUE54(M1_INITCFG1ENABLE),
	.ARGVALUE55(M1_INITCFG2ENABLE),
	.ARGVALUE56(M1_INITCFG3ENABLE),
	.ARGVALUE57(M1_INITCFG4ENABLE),
	.ARGVALUE58(M1_INITCFG5ENABLE),
	.ARGVALUE59(M1_INITCFG6ENABLE),
	.ARGVALUE60(M1_INITCFG7ENABLE),
	.ARGVALUE61(M1_INITCFG8ENABLE),
	.ARGVALUE62(M1_INITCFG9ENABLE),
	.ARGVALUE63(M1_INITCFG10ENABLE),
	.ARGVALUE64(M1_INITCFG11ENABLE),
	.ARGVALUE65(M1_INITCFG12ENABLE),
	.ARGVALUE66(M1_INITCFG13ENABLE),
	.ARGVALUE67(M1_INITCFG14ENABLE),
	.ARGVALUE68(M1_INITCFG15ENABLE)
) master0 (
	// Inputs
	.SYSCLK(SYSCLK),
	.SYSRSTN(SYSRSTN),
	.HREADY(HREADY_M0),
	.HRESP(HRESP_M0[0]),
	.HRDATA(HRDATA_M0),
	// Outputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	.HTRANS(HTRANS_M0),
	.HBURST(),
	.HSEL(),
	.HPROT(),
	.HSIZE(HSIZE_M0),
	.HWRITE(HWRITE_M0),
	.HMASTLOCK(HMASTLOCK_M0),
	.HADDR(HADDR_M0),
	.HWDATA(HWDATA_M0),
	.INTERRUPT(256'b0),
	.GP_OUT(GP_OUT_M0),
	.GP_IN(GP_IN),
	.EXT_WR(),
	.EXT_RD(),
	.EXT_ADDR(),
	.EXT_DATA(),
	.EXT_WAIT(1'b0),
	.FINISHED(FINISHED_master0),
	.FAILED()
);

// control remap signals from master 0 BFM
assign REMAP_M0			= GP_OUT_M0[0];

// signals for testbench request/acknowledgement between masters
assign M0_REQ			= GP_OUT_M0[16];
assign M0_ACK			= GP_OUT_M0[17];


// master 1 BFM
BFM_AHBL  #(
	.VECTFILE(MASTER1_VECTFILE),
	// passing testbench parameters to BFM ARGVALUE* parameters
	.ARGVALUE0(FAMILY),
	.ARGVALUE1(MODE_CFG),
	.ARGVALUE2(M0_AHBSLOT0ENABLE),
	.ARGVALUE3(M0_AHBSLOT1ENABLE),
	.ARGVALUE4(M0_AHBSLOT2ENABLE),
	.ARGVALUE5(M0_AHBSLOT3ENABLE),
	.ARGVALUE6(M0_AHBSLOT4ENABLE),
	.ARGVALUE7(M0_AHBSLOT5ENABLE),
	.ARGVALUE8(M0_AHBSLOT6ENABLE),
	.ARGVALUE9(M0_AHBSLOT7ENABLE),
	.ARGVALUE10(M0_AHBSLOT8ENABLE),
	.ARGVALUE11(M0_AHBSLOT9ENABLE),
	.ARGVALUE12(M0_AHBSLOT10ENABLE),
	.ARGVALUE13(M0_AHBSLOT11ENABLE),
	.ARGVALUE14(M0_AHBSLOT12ENABLE),
	.ARGVALUE15(M0_AHBSLOT13ENABLE),
	.ARGVALUE16(M0_AHBSLOT14ENABLE),
	.ARGVALUE17(M0_AHBSLOT15ENABLE),
	.ARGVALUE18(M1_AHBSLOT0ENABLE),
	.ARGVALUE19(M1_AHBSLOT1ENABLE),
	.ARGVALUE20(M1_AHBSLOT2ENABLE),
	.ARGVALUE21(M1_AHBSLOT3ENABLE),
	.ARGVALUE22(M1_AHBSLOT4ENABLE),
	.ARGVALUE23(M1_AHBSLOT5ENABLE),
	.ARGVALUE24(M1_AHBSLOT6ENABLE),
	.ARGVALUE25(M1_AHBSLOT7ENABLE),
	.ARGVALUE26(M1_AHBSLOT8ENABLE),
	.ARGVALUE27(M1_AHBSLOT9ENABLE),
	.ARGVALUE28(M1_AHBSLOT10ENABLE),
	.ARGVALUE29(M1_AHBSLOT11ENABLE),
	.ARGVALUE30(M1_AHBSLOT12ENABLE),
	.ARGVALUE31(M1_AHBSLOT13ENABLE),
	.ARGVALUE32(M1_AHBSLOT14ENABLE),
	.ARGVALUE33(M1_AHBSLOT15ENABLE),
	.ARGVALUE34(M0_HUGESLOTENABLE),
	.ARGVALUE35(M1_HUGESLOTENABLE),
	.ARGVALUE36(HADDR_SHG_CFG),
	.ARGVALUE37(M0_INITCFG0ENABLE),
	.ARGVALUE38(M0_INITCFG1ENABLE),
	.ARGVALUE39(M0_INITCFG2ENABLE),
	.ARGVALUE40(M0_INITCFG3ENABLE),
	.ARGVALUE41(M0_INITCFG4ENABLE),
	.ARGVALUE42(M0_INITCFG5ENABLE),
	.ARGVALUE43(M0_INITCFG6ENABLE),
	.ARGVALUE44(M0_INITCFG7ENABLE),
	.ARGVALUE45(M0_INITCFG8ENABLE),
	.ARGVALUE46(M0_INITCFG9ENABLE),
	.ARGVALUE47(M0_INITCFG10ENABLE),
	.ARGVALUE48(M0_INITCFG11ENABLE),
	.ARGVALUE49(M0_INITCFG12ENABLE),
	.ARGVALUE50(M0_INITCFG13ENABLE),
	.ARGVALUE51(M0_INITCFG14ENABLE),
	.ARGVALUE52(M0_INITCFG15ENABLE),
	.ARGVALUE53(M1_INITCFG0ENABLE),
	.ARGVALUE54(M1_INITCFG1ENABLE),
	.ARGVALUE55(M1_INITCFG2ENABLE),
	.ARGVALUE56(M1_INITCFG3ENABLE),
	.ARGVALUE57(M1_INITCFG4ENABLE),
	.ARGVALUE58(M1_INITCFG5ENABLE),
	.ARGVALUE59(M1_INITCFG6ENABLE),
	.ARGVALUE60(M1_INITCFG7ENABLE),
	.ARGVALUE61(M1_INITCFG8ENABLE),
	.ARGVALUE62(M1_INITCFG9ENABLE),
	.ARGVALUE63(M1_INITCFG10ENABLE),
	.ARGVALUE64(M1_INITCFG11ENABLE),
	.ARGVALUE65(M1_INITCFG12ENABLE),
	.ARGVALUE66(M1_INITCFG13ENABLE),
	.ARGVALUE67(M1_INITCFG14ENABLE),
	.ARGVALUE68(M1_INITCFG15ENABLE)
) master1 (
	// Inputs
	.SYSCLK(SYSCLK),
	.SYSRSTN(SYSRSTN),
	.HREADY(HREADY_M1),
	.HRESP(HRESP_M1[0]),
	.HRDATA(HRDATA_M1),
	// Outputs
	// using master 0 HCLK,HRESETN to drive slaves & DUT
	//.HCLK(HCLK),
	//.HRESETN(HRESETN),
	.HCLK(),
	.HRESETN(),
	.HTRANS(HTRANS_M1),
	.HBURST(),
	.HSEL(),
	.HPROT(),
	.HSIZE(HSIZE_M1),
	.HWRITE(HWRITE_M1),
	.HMASTLOCK(HMASTLOCK_M1),
	.HADDR(HADDR_M1),
	.HWDATA(HWDATA_M1),
	.INTERRUPT(256'b0),
	.GP_OUT(GP_OUT_M1),
	.GP_IN(GP_IN),
	.EXT_WR(),
	.EXT_RD(),
	.EXT_ADDR(),
	.EXT_DATA(),
	.EXT_WAIT(1'b0),
	.FINISHED(FINISHED_master1),
	.FAILED()
);

// signals for testbench request/acknowledgement between masters
assign M1_REQ			= GP_OUT_M1[18];
assign M1_ACK			= GP_OUT_M1[19];


    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave0 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S0),
	.HSIZE(HSIZE_S0),
	.HTRANS(HTRANS_S0),
	.HWDATA(HWDATA_S0),
	.HREADYIN(HREADYIN_S0),
	.HSEL(HSEL_S0),
	.HADDR(HADDR_S0[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S0),
	.HPROT(HPROT_S0),
	// Output
	.HRDATA(HRDATA_S0),
	.HRESP(HRESP_S0[0]),
	.HREADYOUT(HREADY_S0)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave1 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S1),
	.HSIZE(HSIZE_S1),
	.HTRANS(HTRANS_S1),
	.HWDATA(HWDATA_S1),
	.HREADYIN(HREADYIN_S1),
	.HSEL(HSEL_S1),
	.HADDR(HADDR_S1[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S1),
	.HPROT(HPROT_S1),
	// Output
	.HRDATA(HRDATA_S1),
	.HRESP(HRESP_S1[0]),
	.HREADYOUT(HREADY_S1)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave2 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S2),
	.HSIZE(HSIZE_S2),
	.HTRANS(HTRANS_S2),
	.HWDATA(HWDATA_S2),
	.HREADYIN(HREADYIN_S2),
	.HSEL(HSEL_S2),
	.HADDR(HADDR_S2[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S2),
	.HPROT(HPROT_S2),
	// Output
	.HRDATA(HRDATA_S2),
	.HRESP(HRESP_S2[0]),
	.HREADYOUT(HREADY_S2)
    );


    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave3 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S3),
	.HSIZE(HSIZE_S3),
	.HTRANS(HTRANS_S3),
	.HWDATA(HWDATA_S3),
	.HREADYIN(HREADYIN_S3),
	.HSEL(HSEL_S3),
	.HADDR(HADDR_S3[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S3),
	.HPROT(HPROT_S3),
	// Output
	.HRDATA(HRDATA_S3),
	.HRESP(HRESP_S3[0]),
	.HREADYOUT(HREADY_S3)
    );


    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave4 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S4),
	.HSIZE(HSIZE_S4),
	.HTRANS(HTRANS_S4),
	.HWDATA(HWDATA_S4),
	.HREADYIN(HREADYIN_S4),
	.HSEL(HSEL_S4),
	.HADDR(HADDR_S4[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S4),
	.HPROT(HPROT_S4),
	// Output
	.HRDATA(HRDATA_S4),
	.HRESP(HRESP_S4[0]),
	.HREADYOUT(HREADY_S4)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave5 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S5),
	.HSIZE(HSIZE_S5),
	.HTRANS(HTRANS_S5),
	.HWDATA(HWDATA_S5),
	.HREADYIN(HREADYIN_S5),
	.HSEL(HSEL_S5),
	.HADDR(HADDR_S5[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S5),
	.HPROT(HPROT_S5),
	// Output
	.HRDATA(HRDATA_S5),
	.HRESP(HRESP_S5[0]),
	.HREADYOUT(HREADY_S5)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave6 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S6),
	.HSIZE(HSIZE_S6),
	.HTRANS(HTRANS_S6),
	.HWDATA(HWDATA_S6),
	.HREADYIN(HREADYIN_S6),
	.HSEL(HSEL_S6),
	.HADDR(HADDR_S6[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S6),
	.HPROT(HPROT_S6),
	// Output
	.HRDATA(HRDATA_S6),
	.HRESP(HRESP_S6[0]),
	.HREADYOUT(HREADY_S6)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave7 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S7),
	.HSIZE(HSIZE_S7),
	.HTRANS(HTRANS_S7),
	.HWDATA(HWDATA_S7),
	.HREADYIN(HREADYIN_S7),
	.HSEL(HSEL_S7),
	.HADDR(HADDR_S7[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S7),
	.HPROT(HPROT_S7),
	// Output
	.HRDATA(HRDATA_S7),
	.HRESP(HRESP_S7[0]),
	.HREADYOUT(HREADY_S7)
    );


    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave8 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S8),
	.HSIZE(HSIZE_S8),
	.HTRANS(HTRANS_S8),
	.HWDATA(HWDATA_S8),
	.HREADYIN(HREADYIN_S8),
	.HSEL(HSEL_S8),
	.HADDR(HADDR_S8[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S8),
	.HPROT(HPROT_S8),
	// Output
	.HRDATA(HRDATA_S8),
	.HRESP(HRESP_S8[0]),
	.HREADYOUT(HREADY_S8)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave9 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S9),
	.HSIZE(HSIZE_S9),
	.HTRANS(HTRANS_S9),
	.HWDATA(HWDATA_S9),
	.HREADYIN(HREADYIN_S9),
	.HSEL(HSEL_S9),
	.HADDR(HADDR_S9[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S9),
	.HPROT(HPROT_S9),
	// Output
	.HRDATA(HRDATA_S9),
	.HRESP(HRESP_S9[0]),
	.HREADYOUT(HREADY_S9)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave10 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S10),
	.HSIZE(HSIZE_S10),
	.HTRANS(HTRANS_S10),
	.HWDATA(HWDATA_S10),
	.HREADYIN(HREADYIN_S10),
	.HSEL(HSEL_S10),
	.HADDR(HADDR_S10[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S10),
	.HPROT(HPROT_S10),
	// Output
	.HRDATA(HRDATA_S10),
	.HRESP(HRESP_S10[0]),
	.HREADYOUT(HREADY_S10)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave11 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S11),
	.HSIZE(HSIZE_S11),
	.HTRANS(HTRANS_S11),
	.HWDATA(HWDATA_S11),
	.HREADYIN(HREADYIN_S11),
	.HSEL(HSEL_S11),
	.HADDR(HADDR_S11[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S11),
	.HPROT(HPROT_S11),
	// Output
	.HRDATA(HRDATA_S11),
	.HRESP(HRESP_S11[0]),
	.HREADYOUT(HREADY_S11)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave12 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S12),
	.HSIZE(HSIZE_S12),
	.HTRANS(HTRANS_S12),
	.HWDATA(HWDATA_S12),
	.HREADYIN(HREADYIN_S12),
	.HSEL(HSEL_S12),
	.HADDR(HADDR_S12[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S12),
	.HPROT(HPROT_S12),
	// Output
	.HRDATA(HRDATA_S12),
	.HRESP(HRESP_S12[0]),
	.HREADYOUT(HREADY_S12)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave13 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S13),
	.HSIZE(HSIZE_S13),
	.HTRANS(HTRANS_S13),
	.HWDATA(HWDATA_S13),
	.HREADYIN(HREADYIN_S13),
	.HSEL(HSEL_S13),
	.HADDR(HADDR_S13[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S13),
	.HPROT(HPROT_S13),
	// Output
	.HRDATA(HRDATA_S13),
	.HRESP(HRESP_S13[0]),
	.HREADYOUT(HREADY_S13)
    );


    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave14 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S14),
	.HSIZE(HSIZE_S14),
	.HTRANS(HTRANS_S14),
	.HWDATA(HWDATA_S14),
	.HREADYIN(HREADYIN_S14),
	.HSEL(HSEL_S14),
	.HADDR(HADDR_S14[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S14),
	.HPROT(HPROT_S14),
	// Output
	.HRDATA(HRDATA_S14),
	.HRESP(HRESP_S14[0]),
	.HREADYOUT(HREADY_S14)
    );

    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave15 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_S15),
	.HSIZE(HSIZE_S15),
	.HTRANS(HTRANS_S15),
	.HWDATA(HWDATA_S15),
	.HREADYIN(HREADYIN_S15),
	.HSEL(HSEL_S15),
	.HADDR(HADDR_S15[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_S15),
	.HPROT(HPROT_S15),
	// Output
	.HRDATA(HRDATA_S15),
	.HRESP(HRESP_S15[0]),
	.HREADYOUT(HREADY_S15)
    );

// may need to make this bigger for 'huge' slave
    BFM_AHBSLAVE #(.AWIDTH   (16),
                   .DEPTH    (65536),
                   .INITFILE (" "),
                   .ID       (1),
                   .ENFUNC   (0),
                   .TPD      (5),
                   .DEBUG    (0) ) 
    slave16 (
	// MP7Bridge interface
	// Inputs
	.HCLK(HCLK),
	.HRESETN(HRESETN),
	// AhbFabric interface
	// Inputs
	.HWRITE(HWRITE_SHG),
	.HSIZE(HSIZE_SHG),
	.HTRANS(HTRANS_SHG),
	.HWDATA(HWDATA_SHG),
	.HREADYIN(HREADYIN_SHG),
	.HSEL(HSEL_SHG),
	.HADDR(HADDR_SHG[15:0]),
	.HMASTLOCK(1'b0),
	.HBURST(HBURST_SHG),
	.HPROT(HPROT_SHG),
	// Output
	.HRDATA(HRDATA_SHG),
	.HRESP(HRESP_SHG[0]),
	.HREADYOUT(HREADY_SHG)
    );


endmodule
