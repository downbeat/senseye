`timescale 1ns/1ns
// Copyright 2007 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED 
// Revision Information:
// SVN Revision Information:
// SVN $Revision:  $
module
CoreGPIO
(
PRESETN
,
PCLK
,
PSEL
,
PENABLE
,
PWRITE
,
PSLVERR
,
PREADY
,
PADDR
,
PWDATA
,
PRDATA
,
INT
,
INT_OR
,
GPIO_IN
,
GPIO_OUT
,
GPIO_OE
)
;
parameter
FAMILY
=
17
;
parameter
IO_NUM
=
32
;
parameter
APB_WIDTH
=
32
;
parameter
[
0
:
0
]
OE_TYPE
=
0
;
parameter
[
0
:
0
]
INT_BUS
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_0
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_1
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_2
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_3
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_4
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_5
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_6
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_7
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_8
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_9
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_10
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_11
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_12
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_13
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_14
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_15
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_16
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_17
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_18
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_19
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_20
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_21
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_22
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_23
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_24
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_25
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_26
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_27
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_28
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_29
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_30
=
0
;
parameter
[
0
:
0
]
FIXED_CONFIG_31
=
0
;
parameter
[
1
:
0
]
IO_TYPE_0
=
0
;
parameter
[
1
:
0
]
IO_TYPE_1
=
0
;
parameter
[
1
:
0
]
IO_TYPE_2
=
0
;
parameter
[
1
:
0
]
IO_TYPE_3
=
0
;
parameter
[
1
:
0
]
IO_TYPE_4
=
0
;
parameter
[
1
:
0
]
IO_TYPE_5
=
0
;
parameter
[
1
:
0
]
IO_TYPE_6
=
0
;
parameter
[
1
:
0
]
IO_TYPE_7
=
0
;
parameter
[
1
:
0
]
IO_TYPE_8
=
0
;
parameter
[
1
:
0
]
IO_TYPE_9
=
0
;
parameter
[
1
:
0
]
IO_TYPE_10
=
0
;
parameter
[
1
:
0
]
IO_TYPE_11
=
0
;
parameter
[
1
:
0
]
IO_TYPE_12
=
0
;
parameter
[
1
:
0
]
IO_TYPE_13
=
0
;
parameter
[
1
:
0
]
IO_TYPE_14
=
0
;
parameter
[
1
:
0
]
IO_TYPE_15
=
0
;
parameter
[
1
:
0
]
IO_TYPE_16
=
0
;
parameter
[
1
:
0
]
IO_TYPE_17
=
0
;
parameter
[
1
:
0
]
IO_TYPE_18
=
0
;
parameter
[
1
:
0
]
IO_TYPE_19
=
0
;
parameter
[
1
:
0
]
IO_TYPE_20
=
0
;
parameter
[
1
:
0
]
IO_TYPE_21
=
0
;
parameter
[
1
:
0
]
IO_TYPE_22
=
0
;
parameter
[
1
:
0
]
IO_TYPE_23
=
0
;
parameter
[
1
:
0
]
IO_TYPE_24
=
0
;
parameter
[
1
:
0
]
IO_TYPE_25
=
0
;
parameter
[
1
:
0
]
IO_TYPE_26
=
0
;
parameter
[
1
:
0
]
IO_TYPE_27
=
0
;
parameter
[
1
:
0
]
IO_TYPE_28
=
0
;
parameter
[
1
:
0
]
IO_TYPE_29
=
0
;
parameter
[
1
:
0
]
IO_TYPE_30
=
0
;
parameter
[
1
:
0
]
IO_TYPE_31
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_0
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_1
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_2
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_3
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_4
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_5
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_6
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_7
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_8
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_9
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_10
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_11
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_12
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_13
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_14
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_15
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_16
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_17
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_18
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_19
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_20
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_21
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_22
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_23
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_24
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_25
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_26
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_27
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_28
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_29
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_30
=
0
;
parameter
[
2
:
0
]
IO_INT_TYPE_31
=
0
;
parameter
[
0
:
0
]
IO_VAL_0
=
0
;
parameter
[
0
:
0
]
IO_VAL_1
=
0
;
parameter
[
0
:
0
]
IO_VAL_2
=
0
;
parameter
[
0
:
0
]
IO_VAL_3
=
0
;
parameter
[
0
:
0
]
IO_VAL_4
=
0
;
parameter
[
0
:
0
]
IO_VAL_5
=
0
;
parameter
[
0
:
0
]
IO_VAL_6
=
0
;
parameter
[
0
:
0
]
IO_VAL_7
=
0
;
parameter
[
0
:
0
]
IO_VAL_8
=
0
;
parameter
[
0
:
0
]
IO_VAL_9
=
0
;
parameter
[
0
:
0
]
IO_VAL_10
=
0
;
parameter
[
0
:
0
]
IO_VAL_11
=
0
;
parameter
[
0
:
0
]
IO_VAL_12
=
0
;
parameter
[
0
:
0
]
IO_VAL_13
=
0
;
parameter
[
0
:
0
]
IO_VAL_14
=
0
;
parameter
[
0
:
0
]
IO_VAL_15
=
0
;
parameter
[
0
:
0
]
IO_VAL_16
=
0
;
parameter
[
0
:
0
]
IO_VAL_17
=
0
;
parameter
[
0
:
0
]
IO_VAL_18
=
0
;
parameter
[
0
:
0
]
IO_VAL_19
=
0
;
parameter
[
0
:
0
]
IO_VAL_20
=
0
;
parameter
[
0
:
0
]
IO_VAL_21
=
0
;
parameter
[
0
:
0
]
IO_VAL_22
=
0
;
parameter
[
0
:
0
]
IO_VAL_23
=
0
;
parameter
[
0
:
0
]
IO_VAL_24
=
0
;
parameter
[
0
:
0
]
IO_VAL_25
=
0
;
parameter
[
0
:
0
]
IO_VAL_26
=
0
;
parameter
[
0
:
0
]
IO_VAL_27
=
0
;
parameter
[
0
:
0
]
IO_VAL_28
=
0
;
parameter
[
0
:
0
]
IO_VAL_29
=
0
;
parameter
[
0
:
0
]
IO_VAL_30
=
0
;
parameter
[
0
:
0
]
IO_VAL_31
=
0
;
input
PRESETN
;
input
PCLK
;
input
PSEL
;
input
PENABLE
;
input
PWRITE
;
output
PSLVERR
;
output
PREADY
;
input
[
7
:
0
]
PADDR
;
input
[
APB_WIDTH
-
1
:
0
]
PWDATA
;
output
[
APB_WIDTH
-
1
:
0
]
PRDATA
;
output
[
IO_NUM
-
1
:
0
]
INT
;
output
INT_OR
;
input
[
IO_NUM
-
1
:
0
]
GPIO_IN
;
output
[
IO_NUM
-
1
:
0
]
GPIO_OUT
;
output
[
IO_NUM
-
1
:
0
]
GPIO_OE
;
parameter
[
0
:
31
]
CGPIOO
=
(
{
FIXED_CONFIG_0
,
FIXED_CONFIG_1
,
FIXED_CONFIG_2
,
FIXED_CONFIG_3
,
FIXED_CONFIG_4
,
FIXED_CONFIG_5
,
FIXED_CONFIG_6
,
FIXED_CONFIG_7
,
FIXED_CONFIG_8
,
FIXED_CONFIG_9
,
FIXED_CONFIG_10
,
FIXED_CONFIG_11
,
FIXED_CONFIG_12
,
FIXED_CONFIG_13
,
FIXED_CONFIG_14
,
FIXED_CONFIG_15
,
FIXED_CONFIG_16
,
FIXED_CONFIG_17
,
FIXED_CONFIG_18
,
FIXED_CONFIG_19
,
FIXED_CONFIG_20
,
FIXED_CONFIG_21
,
FIXED_CONFIG_22
,
FIXED_CONFIG_23
,
FIXED_CONFIG_24
,
FIXED_CONFIG_25
,
FIXED_CONFIG_26
,
FIXED_CONFIG_27
,
FIXED_CONFIG_28
,
FIXED_CONFIG_29
,
FIXED_CONFIG_30
,
FIXED_CONFIG_31
}
)
;
parameter
[
0
:
95
]
CGPIOI
=
(
{
IO_INT_TYPE_0
,
IO_INT_TYPE_1
,
IO_INT_TYPE_2
,
IO_INT_TYPE_3
,
IO_INT_TYPE_4
,
IO_INT_TYPE_5
,
IO_INT_TYPE_6
,
IO_INT_TYPE_7
,
IO_INT_TYPE_8
,
IO_INT_TYPE_9
,
IO_INT_TYPE_10
,
IO_INT_TYPE_11
,
IO_INT_TYPE_12
,
IO_INT_TYPE_13
,
IO_INT_TYPE_14
,
IO_INT_TYPE_15
,
IO_INT_TYPE_16
,
IO_INT_TYPE_17
,
IO_INT_TYPE_18
,
IO_INT_TYPE_19
,
IO_INT_TYPE_20
,
IO_INT_TYPE_21
,
IO_INT_TYPE_22
,
IO_INT_TYPE_23
,
IO_INT_TYPE_24
,
IO_INT_TYPE_25
,
IO_INT_TYPE_26
,
IO_INT_TYPE_27
,
IO_INT_TYPE_28
,
IO_INT_TYPE_29
,
IO_INT_TYPE_30
,
IO_INT_TYPE_31
}
)
;
parameter
[
0
:
63
]
CGPIOl
=
(
{
IO_TYPE_0
,
IO_TYPE_1
,
IO_TYPE_2
,
IO_TYPE_3
,
IO_TYPE_4
,
IO_TYPE_5
,
IO_TYPE_6
,
IO_TYPE_7
,
IO_TYPE_8
,
IO_TYPE_9
,
IO_TYPE_10
,
IO_TYPE_11
,
IO_TYPE_12
,
IO_TYPE_13
,
IO_TYPE_14
,
IO_TYPE_15
,
IO_TYPE_16
,
IO_TYPE_17
,
IO_TYPE_18
,
IO_TYPE_19
,
IO_TYPE_20
,
IO_TYPE_21
,
IO_TYPE_22
,
IO_TYPE_23
,
IO_TYPE_24
,
IO_TYPE_25
,
IO_TYPE_26
,
IO_TYPE_27
,
IO_TYPE_28
,
IO_TYPE_29
,
IO_TYPE_30
,
IO_TYPE_31
}
)
;
parameter
[
0
:
31
]
CGPIOOI
=
(
{
IO_VAL_0
,
IO_VAL_1
,
IO_VAL_2
,
IO_VAL_3
,
IO_VAL_4
,
IO_VAL_5
,
IO_VAL_6
,
IO_VAL_7
,
IO_VAL_8
,
IO_VAL_9
,
IO_VAL_10
,
IO_VAL_11
,
IO_VAL_12
,
IO_VAL_13
,
IO_VAL_14
,
IO_VAL_15
,
IO_VAL_16
,
IO_VAL_17
,
IO_VAL_18
,
IO_VAL_19
,
IO_VAL_20
,
IO_VAL_21
,
IO_VAL_22
,
IO_VAL_23
,
IO_VAL_24
,
IO_VAL_25
,
IO_VAL_26
,
IO_VAL_27
,
IO_VAL_28
,
IO_VAL_29
,
IO_VAL_30
,
IO_VAL_31
}
)
;
reg
[
7
:
0
]
CGPIOII
[
0
:
IO_NUM
-
1
]
;
reg
[
31
:
0
]
CGPIOlI
;
reg
[
32
-
1
:
0
]
CGPIOOl
;
reg
[
32
-
1
:
0
]
CGPIOIl
;
wire
[
32
-
1
:
0
]
CGPIOll
;
wire
[
IO_NUM
-
1
:
0
]
CGPIOO0
;
wire
[
IO_NUM
-
1
:
0
]
CGPIOI0
;
wire
[
APB_WIDTH
-
1
:
0
]
CGPIOl0
;
reg
[
IO_NUM
-
1
:
0
]
CGPIOO1
;
reg
[
IO_NUM
-
1
:
0
]
CGPIOI1
;
reg
[
IO_NUM
-
1
:
0
]
CGPIOl1
;
reg
[
IO_NUM
-
1
:
0
]
CGPIOOOI
;
reg
[
IO_NUM
-
1
:
0
]
CGPIOIOI
;
reg
[
IO_NUM
-
1
:
0
]
CGPIOlOI
;
wire
[
IO_NUM
-
1
:
0
]
CGPIOOII
;
wire
[
IO_NUM
-
1
:
0
]
CGPIOIII
;
wire
[
IO_NUM
-
1
:
0
]
CGPIOlII
;
wire
[
IO_NUM
-
1
:
0
]
CGPIOOlI
;
wire
[
IO_NUM
-
1
:
0
]
CGPIOIlI
;
wire
[
31
:
0
]
CGPIOllI
;
wire
[
5
:
0
]
CGPIOO0I
;
wire
CGPIOI0I
;
wire
[
7
:
0
]
CGPIOl0I
;
assign
CGPIOI0I
=
1
'b
0
;
assign
CGPIOl0I
=
8
'h
00
;
assign
PSLVERR
=
1
'b
0
;
assign
PREADY
=
1
'b
1
;
assign
PRDATA
[
APB_WIDTH
-
1
:
0
]
=
CGPIOl0
[
APB_WIDTH
-
1
:
0
]
;
generate
if
(
INT_BUS
==
1
)
assign
INT_OR
=
|
CGPIOOlI
;
else
assign
INT_OR
=
1
'b
0
;
endgenerate
generate
if
(
IO_NUM
<
32
)
begin
:
CGPIOO1I
genvar
J
;
for
(
J
=
IO_NUM
;
J
<=
31
;
J
=
J
+
1
)
begin
:
CGPIOI1I
assign
CGPIOll
[
J
]
=
1
'b
0
;
always
@
*
begin
CGPIOIl
[
J
]
<=
CGPIOI0I
;
CGPIOOl
[
J
]
<=
CGPIOI0I
;
end
end
end
endgenerate
generate
begin
:
CGPIOl1I
genvar
CGPIOOOl
;
for
(
CGPIOOOl
=
0
;
CGPIOOOl
<=
(
IO_NUM
-
1
)
;
CGPIOOOl
=
CGPIOOOl
+
1
)
begin
:
CGPIOIOl
assign
CGPIOOII
[
CGPIOOOl
]
=
CGPIOI1
[
CGPIOOOl
]
;
assign
CGPIOlII
[
CGPIOOOl
]
=
CGPIOl1
[
CGPIOOOl
]
;
assign
CGPIOIII
[
CGPIOOOl
]
=
(
~
CGPIOl1
[
CGPIOOOl
]
)
;
assign
INT
[
CGPIOOOl
]
=
CGPIOOlI
[
CGPIOOOl
]
;
assign
GPIO_OE
=
CGPIOI0
;
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
begin
CGPIOO1
[
CGPIOOOl
]
<=
1
'b
0
;
CGPIOI1
[
CGPIOOOl
]
<=
1
'b
0
;
end
else
begin
CGPIOO1
[
CGPIOOOl
]
<=
GPIO_IN
[
CGPIOOOl
]
;
CGPIOI1
[
CGPIOOOl
]
<=
CGPIOO1
[
CGPIOOOl
]
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOl1
[
CGPIOOOl
]
<=
1
'b
0
;
else
CGPIOl1
[
CGPIOOOl
]
<=
CGPIOOII
[
CGPIOOOl
]
;
if
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
begin
:
CGPIOlOl
assign
CGPIOIlI
[
CGPIOOOl
]
=
(
(
CGPIOII
[
CGPIOOOl
]
[
7
:
5
]
==
3
'b
000
)
)
?
CGPIOlII
[
CGPIOOOl
]
:
(
(
CGPIOII
[
CGPIOOOl
]
[
7
:
5
]
==
3
'b
001
)
)
?
CGPIOIII
[
CGPIOOOl
]
:
(
(
CGPIOII
[
CGPIOOOl
]
[
7
:
5
]
==
3
'b
010
)
)
?
CGPIOOOI
[
CGPIOOOl
]
:
(
(
CGPIOII
[
CGPIOOOl
]
[
7
:
5
]
==
3
'b
011
)
)
?
CGPIOlOI
[
CGPIOOOl
]
:
(
(
CGPIOII
[
CGPIOOOl
]
[
7
:
5
]
==
3
'b
100
)
)
?
CGPIOIOI
[
CGPIOOOl
]
:
1
'b
0
;
assign
CGPIOOlI
[
CGPIOOOl
]
=
(
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
?
CGPIOIlI
[
CGPIOOOl
]
:
1
'b
0
;
end
if
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
begin
:
CGPIOOIl
assign
CGPIOIlI
[
CGPIOOOl
]
=
(
(
CGPIOI
[
3
*
CGPIOOOl
:
3
*
CGPIOOOl
+
2
]
==
3
'b
000
)
)
?
CGPIOlII
[
CGPIOOOl
]
:
(
(
CGPIOI
[
3
*
CGPIOOOl
:
3
*
CGPIOOOl
+
2
]
==
3
'b
001
)
)
?
CGPIOIII
[
CGPIOOOl
]
:
(
(
CGPIOI
[
3
*
CGPIOOOl
:
3
*
CGPIOOOl
+
2
]
==
3
'b
010
)
)
?
CGPIOOOI
[
CGPIOOOl
]
:
(
(
CGPIOI
[
3
*
CGPIOOOl
:
3
*
CGPIOOOl
+
2
]
==
3
'b
011
)
)
?
CGPIOlOI
[
CGPIOOOl
]
:
(
(
CGPIOI
[
3
*
CGPIOOOl
:
3
*
CGPIOOOl
+
2
]
==
3
'b
100
)
)
?
CGPIOIOI
[
CGPIOOOl
]
:
1
'b
0
;
assign
CGPIOOlI
[
CGPIOOOl
]
=
(
(
CGPIOI
[
3
*
CGPIOOOl
:
3
*
CGPIOOOl
+
2
]
!=
3
'b
111
)
)
?
CGPIOIlI
[
CGPIOOOl
]
:
1
'b
0
;
end
if
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
begin
:
CGPIOIIl
assign
CGPIOll
[
CGPIOOOl
]
=
(
(
CGPIOII
[
CGPIOOOl
]
[
1
]
==
1
'b
1
)
)
?
CGPIOl1
[
CGPIOOOl
]
:
1
'b
0
;
end
if
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
begin
:
CGPIOlIl
assign
CGPIOll
[
CGPIOOOl
]
=
(
(
CGPIOl
[
2
*
CGPIOOOl
:
2
*
CGPIOOOl
+
1
]
!=
2
'b
01
)
)
?
CGPIOl1
[
CGPIOOOl
]
:
1
'b
0
;
end
if
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
begin
:
CGPIOOll
assign
CGPIOO0
[
CGPIOOOl
]
=
(
(
CGPIOII
[
CGPIOOOl
]
[
0
]
==
1
'b
1
)
)
?
CGPIOIl
[
CGPIOOOl
]
:
1
'b
0
;
assign
CGPIOI0
[
CGPIOOOl
]
=
(
(
CGPIOII
[
CGPIOOOl
]
[
2
]
==
1
'b
1
)
&&
(
CGPIOII
[
CGPIOOOl
]
[
0
]
==
1
'b
1
)
)
?
1
'b
1
:
1
'b
0
;
end
if
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
begin
:
CGPIOIll
assign
CGPIOO0
[
CGPIOOOl
]
=
(
(
CGPIOl
[
2
*
CGPIOOOl
:
2
*
CGPIOOOl
+
1
]
!=
2
'b
00
)
)
?
CGPIOIl
[
CGPIOOOl
]
:
1
'b
0
;
assign
CGPIOI0
[
CGPIOOOl
]
=
1
'b
1
;
end
if
(
OE_TYPE
==
0
)
begin
:
CGPIOlll
assign
GPIO_OUT
[
CGPIOOOl
]
=
CGPIOO0
[
CGPIOOOl
]
;
end
if
(
OE_TYPE
==
1
)
begin
:
CGPIOO0l
assign
GPIO_OUT
[
CGPIOOOl
]
=
(
(
CGPIOI0
[
CGPIOOOl
]
==
1
'b
1
)
)
?
CGPIOO0
[
CGPIOOOl
]
:
1
'b
Z
;
end
if
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
begin
:
CGPIOI0l
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
begin
if
(
PRESETN
==
1
'b
0
)
CGPIOII
[
CGPIOOOl
]
[
7
:
0
]
<=
8
'h
00
;
else
begin
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
2
]
==
CGPIOOOl
)
)
CGPIOII
[
CGPIOOOl
]
[
7
:
0
]
<=
PWDATA
[
7
:
0
]
;
else
CGPIOII
[
CGPIOOOl
]
[
7
:
0
]
<=
CGPIOII
[
CGPIOOOl
]
[
7
:
0
]
;
end
end
end
else
begin
always
@
*
begin
CGPIOII
[
CGPIOOOl
]
[
7
:
0
]
<=
CGPIOl0I
;
end
end
if
(
APB_WIDTH
==
32
)
begin
:
CGPIOl0l
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOOOI
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
&
(
CGPIOI
[
(
3
*
CGPIOOOl
)
:
(
3
*
CGPIOOOl
+
2
)
]
==
3
'b
010
)
)
|
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
&
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
)
begin
if
(
(
CGPIOOII
[
CGPIOOOl
]
==
1
'b
1
)
&
(
(
~
CGPIOl1
[
CGPIOOOl
]
)
==
1
'b
1
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
1
'b
1
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
;
end
else
CGPIOOOI
[
CGPIOOOl
]
<=
1
'b
0
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOlOI
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
&
(
CGPIOI
[
(
3
*
CGPIOOOl
)
:
(
3
*
CGPIOOOl
+
2
)
]
==
3
'b
011
)
)
|
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
&
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
)
begin
if
(
(
(
~
CGPIOOII
[
CGPIOOOl
]
)
==
1
'b
1
)
&
(
CGPIOl1
[
CGPIOOOl
]
==
1
'b
1
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
1
'b
1
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
;
end
else
CGPIOlOI
[
CGPIOOOl
]
<=
1
'b
0
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOIOI
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
&
(
CGPIOI
[
(
3
*
CGPIOOOl
)
:
(
3
*
CGPIOOOl
+
2
)
]
==
3
'b
100
)
)
|
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
&
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
)
begin
if
(
(
CGPIOOII
[
CGPIOOOl
]
==
1
'b
1
)
^
(
CGPIOl1
[
CGPIOOOl
]
==
1
'b
1
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
1
'b
1
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
;
end
else
CGPIOIOI
[
CGPIOOOl
]
<=
1
'b
0
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOOl
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
)
case
(
PADDR
[
7
:
0
]
)
8
'h
80
:
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOl
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
default
:
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOlI
[
CGPIOOOl
]
;
endcase
else
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOlI
[
CGPIOOOl
]
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOIl
[
CGPIOOOl
]
<=
CGPIOOI
[
CGPIOOOl
]
;
else
begin
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
)
case
(
PADDR
[
7
:
0
]
)
8
'h
A0
:
CGPIOIl
[
CGPIOOOl
]
<=
PWDATA
[
CGPIOOOl
]
;
default
:
CGPIOIl
[
CGPIOOOl
]
<=
CGPIOIl
[
CGPIOOOl
]
;
endcase
else
CGPIOIl
[
CGPIOOOl
]
<=
CGPIOIl
[
CGPIOOOl
]
;
end
end
if
(
APB_WIDTH
==
16
)
begin
:
CGPIOO1l
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOOOI
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
&
(
CGPIOI
[
(
3
*
CGPIOOOl
)
:
(
3
*
CGPIOOOl
+
2
)
]
==
3
'b
010
)
)
|
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
&
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
)
begin
if
(
(
CGPIOOII
[
CGPIOOOl
]
==
1
'b
1
)
&
(
(
~
CGPIOl1
[
CGPIOOOl
]
)
==
1
'b
1
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
1
'b
1
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
&
(
CGPIOOOl
<
16
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
84
)
&
(
CGPIOOOl
>=
16
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
16
]
)
)
;
else
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
;
end
else
CGPIOOOI
[
CGPIOOOl
]
<=
1
'b
0
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOlOI
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
&
(
CGPIOI
[
(
3
*
CGPIOOOl
)
:
(
3
*
CGPIOOOl
+
2
)
]
==
3
'b
011
)
)
|
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
&
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
)
begin
if
(
(
(
~
CGPIOOII
[
CGPIOOOl
]
)
==
1
'b
1
)
&
(
CGPIOl1
[
CGPIOOOl
]
==
1
'b
1
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
1
'b
1
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
&
(
CGPIOOOl
<
16
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
84
)
&
(
CGPIOOOl
>=
16
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
16
]
)
)
;
else
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
;
end
else
CGPIOlOI
[
CGPIOOOl
]
<=
1
'b
0
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOIOI
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
&
(
CGPIOI
[
(
3
*
CGPIOOOl
)
:
(
3
*
CGPIOOOl
+
2
)
]
==
3
'b
100
)
)
|
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
&
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
)
begin
if
(
(
CGPIOOII
[
CGPIOOOl
]
==
1
'b
1
)
^
(
CGPIOl1
[
CGPIOOOl
]
==
1
'b
1
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
1
'b
1
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
&
(
CGPIOOOl
<
16
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
84
)
&
(
CGPIOOOl
>=
16
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
16
]
)
)
;
else
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
;
end
else
CGPIOIOI
[
CGPIOOOl
]
<=
1
'b
0
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOOl
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
&
(
CGPIOOOl
<
16
)
)
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOl
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
84
)
&
(
CGPIOOOl
>=
16
)
)
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOl
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
16
]
)
)
;
else
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOlI
[
CGPIOOOl
]
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOIl
[
CGPIOOOl
]
<=
CGPIOOI
[
CGPIOOOl
]
;
else
begin
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
A0
)
&
(
CGPIOOOl
<
16
)
)
CGPIOIl
[
CGPIOOOl
]
<=
PWDATA
[
CGPIOOOl
]
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
A4
)
&
(
CGPIOOOl
>=
16
)
)
CGPIOIl
[
CGPIOOOl
]
<=
PWDATA
[
CGPIOOOl
-
16
]
;
else
CGPIOIl
[
CGPIOOOl
]
<=
CGPIOIl
[
CGPIOOOl
]
;
end
end
if
(
APB_WIDTH
==
8
)
begin
:
CGPIOI1l
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOOOI
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
&
(
CGPIOI
[
(
3
*
CGPIOOOl
)
:
(
3
*
CGPIOOOl
+
2
)
]
==
3
'b
010
)
)
|
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
&
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
)
begin
if
(
(
CGPIOOII
[
CGPIOOOl
]
==
1
'b
1
)
&
(
(
~
CGPIOl1
[
CGPIOOOl
]
)
==
1
'b
1
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
1
'b
1
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
&
(
CGPIOOOl
<
8
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
84
)
&
(
CGPIOOOl
>=
8
)
&
(
CGPIOOOl
<
16
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
8
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
88
)
&
(
CGPIOOOl
>=
16
)
&
(
CGPIOOOl
<
24
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
16
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
8C
)
&
(
CGPIOOOl
>=
24
)
)
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
24
]
)
)
;
else
CGPIOOOI
[
CGPIOOOl
]
<=
CGPIOOOI
[
CGPIOOOl
]
;
end
else
CGPIOOOI
[
CGPIOOOl
]
<=
1
'b
0
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOlOI
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
&
(
CGPIOI
[
(
3
*
CGPIOOOl
)
:
(
3
*
CGPIOOOl
+
2
)
]
==
3
'b
011
)
)
|
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
&
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
)
begin
if
(
(
(
~
CGPIOOII
[
CGPIOOOl
]
)
==
1
'b
1
)
&
(
CGPIOl1
[
CGPIOOOl
]
==
1
'b
1
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
1
'b
1
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
&
(
CGPIOOOl
<
8
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
84
)
&
(
CGPIOOOl
>=
8
)
&
(
CGPIOOOl
<
16
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
8
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
88
)
&
(
CGPIOOOl
>=
16
)
&
(
CGPIOOOl
<
24
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
16
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
8C
)
&
(
CGPIOOOl
>=
24
)
)
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
24
]
)
)
;
else
CGPIOlOI
[
CGPIOOOl
]
<=
CGPIOlOI
[
CGPIOOOl
]
;
end
else
CGPIOlOI
[
CGPIOOOl
]
<=
1
'b
0
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOIOI
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
1
)
&
(
CGPIOI
[
(
3
*
CGPIOOOl
)
:
(
3
*
CGPIOOOl
+
2
)
]
==
3
'b
100
)
)
|
(
(
CGPIOO
[
CGPIOOOl
]
==
1
'b
0
)
&
(
CGPIOII
[
CGPIOOOl
]
[
3
]
==
1
'b
1
)
)
)
begin
if
(
(
CGPIOOII
[
CGPIOOOl
]
==
1
'b
1
)
^
(
CGPIOl1
[
CGPIOOOl
]
==
1
'b
1
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
1
'b
1
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
&
(
CGPIOOOl
<
8
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
84
)
&
(
CGPIOOOl
>=
8
)
&
(
CGPIOOOl
<
16
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
8
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
88
)
&
(
CGPIOOOl
>=
16
)
&
(
CGPIOOOl
<
24
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
16
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
8C
)
&
(
CGPIOOOl
>=
24
)
)
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
24
]
)
)
;
else
CGPIOIOI
[
CGPIOOOl
]
<=
CGPIOIOI
[
CGPIOOOl
]
;
end
else
CGPIOIOI
[
CGPIOOOl
]
<=
1
'b
0
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOOl
[
CGPIOOOl
]
<=
1
'b
0
;
else
begin
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
80
)
&
(
CGPIOOOl
<
8
)
)
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOl
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
84
)
&
(
CGPIOOOl
>=
8
)
&
(
CGPIOOOl
<
16
)
)
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOl
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
8
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
88
)
&
(
CGPIOOOl
>=
16
)
&
(
CGPIOOOl
<
24
)
)
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOl
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
16
]
)
)
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
8C
)
&
(
CGPIOOOl
>=
24
)
)
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOl
[
CGPIOOOl
]
&
(
(
~
PWDATA
[
CGPIOOOl
-
24
]
)
)
;
else
CGPIOOl
[
CGPIOOOl
]
<=
CGPIOOlI
[
CGPIOOOl
]
;
end
always
@
(
posedge
PCLK
or
negedge
PRESETN
)
if
(
PRESETN
==
1
'b
0
)
CGPIOIl
[
CGPIOOOl
]
<=
CGPIOOI
[
CGPIOOOl
]
;
else
begin
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
A0
)
&
(
CGPIOOOl
<
8
)
)
CGPIOIl
[
CGPIOOOl
]
<=
PWDATA
[
CGPIOOOl
]
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
A4
)
&
(
CGPIOOOl
>=
8
)
&
(
CGPIOOOl
<
16
)
)
CGPIOIl
[
CGPIOOOl
]
<=
PWDATA
[
CGPIOOOl
-
8
]
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
A8
)
&
(
CGPIOOOl
>=
16
)
&
(
CGPIOOOl
<
24
)
)
CGPIOIl
[
CGPIOOOl
]
<=
PWDATA
[
CGPIOOOl
-
16
]
;
else
if
(
(
PSEL
==
1
'b
1
)
&
(
PWRITE
==
1
'b
1
)
&
(
PENABLE
==
1
'b
1
)
&
(
PADDR
[
7
:
0
]
==
8
'h
AC
)
&
(
CGPIOOOl
>=
24
)
)
CGPIOIl
[
CGPIOOOl
]
<=
PWDATA
[
CGPIOOOl
-
24
]
;
else
CGPIOIl
[
CGPIOOOl
]
<=
CGPIOIl
[
CGPIOOOl
]
;
end
end
end
end
endgenerate
assign
CGPIOO0I
[
5
:
0
]
=
PADDR
[
7
:
2
]
;
assign
CGPIOllI
=
CGPIOO0I
;
always
@
*
case
(
CGPIOllI
)
0
,
1
,
2
,
3
,
4
,
5
,
6
,
7
,
8
,
9
,
10
,
11
,
12
,
13
,
14
,
15
,
16
,
17
,
18
,
19
,
20
,
21
,
22
,
23
,
24
,
25
,
26
,
27
,
28
,
29
,
30
,
31
:
CGPIOlI
[
31
:
0
]
<=
{
1
'b
0
,
CGPIOII
[
CGPIOllI
]
[
7
:
0
]
}
;
default
:
CGPIOlI
[
31
:
0
]
<=
{
32
{
1
'b
0
}
}
;
endcase
generate
if
(
APB_WIDTH
==
32
)
begin
:
CGPIOl1l
assign
CGPIOl0
[
31
:
0
]
=
(
(
PADDR
[
7
:
0
]
<
8
'h
80
)
)
?
CGPIOlI
[
31
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
80
)
)
?
CGPIOOl
[
31
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
90
)
)
?
CGPIOll
[
31
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
A0
)
)
?
CGPIOIl
[
31
:
0
]
:
32
'h
00000000
;
end
endgenerate
generate
if
(
APB_WIDTH
==
16
)
begin
:
CGPIOOO0
assign
CGPIOl0
[
15
:
0
]
=
(
(
PADDR
[
7
:
0
]
<
8
'h
80
)
)
?
CGPIOlI
[
15
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
80
)
)
?
CGPIOOl
[
15
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
84
)
)
?
CGPIOOl
[
31
:
16
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
90
)
)
?
CGPIOll
[
15
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
94
)
)
?
CGPIOll
[
31
:
16
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
A0
)
)
?
CGPIOIl
[
15
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
A4
)
)
?
CGPIOIl
[
31
:
16
]
:
16
'h
0000
;
end
endgenerate
generate
if
(
APB_WIDTH
==
8
)
begin
:
CGPIOIO0
assign
CGPIOl0
[
7
:
0
]
=
(
(
PADDR
[
7
:
0
]
<
8
'h
80
)
)
?
CGPIOlI
[
7
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
80
)
)
?
CGPIOOl
[
7
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
84
)
)
?
CGPIOOl
[
15
:
8
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
88
)
)
?
CGPIOOl
[
23
:
16
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
8C
)
)
?
CGPIOOl
[
31
:
24
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
90
)
)
?
CGPIOll
[
7
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
94
)
)
?
CGPIOll
[
15
:
8
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
98
)
)
?
CGPIOll
[
23
:
16
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
9C
)
)
?
CGPIOll
[
31
:
24
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
A0
)
)
?
CGPIOIl
[
7
:
0
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
A4
)
)
?
CGPIOIl
[
15
:
8
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
A8
)
)
?
CGPIOIl
[
23
:
16
]
:
(
(
PADDR
[
7
:
0
]
==
8
'h
AC
)
)
?
CGPIOIl
[
31
:
24
]
:
8
'h
00
;
end
endgenerate
endmodule
