`timescale 1ns/1ps
module
CoreInterrupt
(
PCLK
,
PRESETn
,
PENABLE
,
PSEL
,
PADDR
,
PWRITE
,
PWDATA
,
PRDATA
,
fiqSource7
,
fiqSource6
,
fiqSource5
,
fiqSource4
,
fiqSource3
,
fiqSource2
,
fiqSource1
,
fiqSource0
,
irqSource31
,
irqSource30
,
irqSource29
,
irqSource28
,
irqSource27
,
irqSource26
,
irqSource25
,
irqSource24
,
irqSource23
,
irqSource22
,
irqSource21
,
irqSource20
,
irqSource19
,
irqSource18
,
irqSource17
,
irqSource16
,
irqSource15
,
irqSource14
,
irqSource13
,
irqSource12
,
irqSource11
,
irqSource10
,
irqSource9
,
irqSource8
,
irqSource7
,
irqSource6
,
irqSource5
,
irqSource4
,
irqSource3
,
irqSource2
,
irqSource1
,
irqSource0
,
IRQ
,
FIQ
)
;
`define CoreInterrupt_O  \
4 \
'h \
0
`define CoreInterrupt_I  \
4 \
'h \
1
`define CoreInterrupt_l  \
4 \
'h \
2
`define CoreInterrupt_OI  \
4 \
'h \
3
`define CoreInterrupt_II  \
4 \
'h \
4
`define CoreInterrupt_lI  \
4 \
'h \
5
`define CoreInterrupt_Ol  \
4 \
'h \
6
`define CoreInterrupt_Il  \
4 \
'h \
7
`define CoreInterrupt_ll  \
4 \
'h \
8
`define CoreInterrupt_O0  \
4 \
'h \
9
`define CoreInterrupt_I0  \
4 \
'h \
a
`define CoreInterrupt_l0  \
4 \
'h \
b
parameter
NUMIRQSRC
=
8
;
parameter
NUMFIQSRC
=
0
;
parameter
IRQPOLARITY
=
0
;
parameter
FIQPOLARITY
=
0
;
input
PCLK
;
input
PRESETn
;
input
PENABLE
;
input
PSEL
;
input
[
5
:
2
]
PADDR
;
input
PWRITE
;
input
[
31
:
0
]
PWDATA
;
output
[
31
:
0
]
PRDATA
;
input
fiqSource7
;
input
fiqSource6
;
input
fiqSource5
;
input
fiqSource4
;
input
fiqSource3
;
input
fiqSource2
;
input
fiqSource1
;
input
fiqSource0
;
input
irqSource31
;
input
irqSource30
;
input
irqSource29
;
input
irqSource28
;
input
irqSource27
;
input
irqSource26
;
input
irqSource25
;
input
irqSource24
;
input
irqSource23
;
input
irqSource22
;
input
irqSource21
;
input
irqSource20
;
input
irqSource19
;
input
irqSource18
;
input
irqSource17
;
input
irqSource16
;
input
irqSource15
;
input
irqSource14
;
input
irqSource13
;
input
irqSource12
;
input
irqSource11
;
input
irqSource10
;
input
irqSource9
;
input
irqSource8
;
input
irqSource7
;
input
irqSource6
;
input
irqSource5
;
input
irqSource4
;
input
irqSource3
;
input
irqSource2
;
input
irqSource1
;
input
irqSource0
;
output
IRQ
;
output
FIQ
;
wire
PCLK
;
wire
PRESETn
;
wire
PENABLE
;
wire
PSEL
;
wire
[
5
:
2
]
PADDR
;
wire
PWRITE
;
wire
[
31
:
0
]
PWDATA
;
wire
[
31
:
0
]
PRDATA
;
wire
[
7
:
0
]
CoreInterrupt_O1
;
wire
[
31
:
0
]
CoreInterrupt_I1
;
wire
IRQ
;
wire
FIQ
;
wire
[
31
:
0
]
CoreInterrupt_l1
;
reg
[
31
:
0
]
CoreInterrupt_OOI
;
wire
CoreInterrupt_IOI
;
reg
[
31
:
0
]
CoreInterrupt_lOI
;
wire
[
7
:
0
]
CoreInterrupt_OII
;
wire
[
31
:
0
]
CoreInterrupt_III
;
wire
CoreInterrupt_lII
;
wire
[
7
:
0
]
CoreInterrupt_OlI
;
wire
[
7
:
0
]
CoreInterrupt_IlI
;
wire
[
7
:
0
]
CoreInterrupt_llI
;
reg
[
7
:
0
]
CoreInterrupt_O0I
;
reg
[
7
:
0
]
CoreInterrupt_I0I
;
wire
[
31
:
0
]
CoreInterrupt_l0I
;
wire
[
31
:
0
]
CoreInterrupt_O1I
;
wire
[
31
:
0
]
CoreInterrupt_I1I
;
reg
[
31
:
0
]
CoreInterrupt_l1I
;
reg
[
31
:
0
]
CoreInterrupt_OOl
;
wire
[
7
:
0
]
CoreInterrupt_IOl
;
wire
[
31
:
0
]
CoreInterrupt_lOl
;
assign
CoreInterrupt_O1
=
{
fiqSource7
,
fiqSource6
,
fiqSource5
,
fiqSource4
,
fiqSource3
,
fiqSource2
,
fiqSource1
,
fiqSource0
}
;
assign
CoreInterrupt_I1
=
{
irqSource31
,
irqSource30
,
irqSource29
,
irqSource28
,
irqSource27
,
irqSource26
,
irqSource25
,
irqSource24
,
irqSource23
,
irqSource22
,
irqSource21
,
irqSource20
,
irqSource19
,
irqSource18
,
irqSource17
,
irqSource16
,
irqSource15
,
irqSource14
,
irqSource13
,
irqSource12
,
irqSource11
,
irqSource10
,
irqSource9
,
irqSource8
,
irqSource7
,
irqSource6
,
irqSource5
,
irqSource4
,
irqSource3
,
irqSource2
,
irqSource1
,
irqSource0
}
;
assign
CoreInterrupt_lII
=
(
PWRITE
&&
PSEL
&&
!
PENABLE
)
;
assign
CoreInterrupt_III
=
(
NUMIRQSRC
==
32
)
?
32
'h
ffffffff
:
(
NUMIRQSRC
==
31
)
?
32
'h
7fffffff
:
(
NUMIRQSRC
==
30
)
?
32
'h
3fffffff
:
(
NUMIRQSRC
==
29
)
?
32
'h
1fffffff
:
(
NUMIRQSRC
==
28
)
?
32
'h
0fffffff
:
(
NUMIRQSRC
==
27
)
?
32
'h
07ffffff
:
(
NUMIRQSRC
==
26
)
?
32
'h
03ffffff
:
(
NUMIRQSRC
==
25
)
?
32
'h
01ffffff
:
(
NUMIRQSRC
==
24
)
?
32
'h
00ffffff
:
(
NUMIRQSRC
==
23
)
?
32
'h
007fffff
:
(
NUMIRQSRC
==
22
)
?
32
'h
003fffff
:
(
NUMIRQSRC
==
21
)
?
32
'h
001fffff
:
(
NUMIRQSRC
==
20
)
?
32
'h
000fffff
:
(
NUMIRQSRC
==
19
)
?
32
'h
0007ffff
:
(
NUMIRQSRC
==
18
)
?
32
'h
0003ffff
:
(
NUMIRQSRC
==
17
)
?
32
'h
0001ffff
:
(
NUMIRQSRC
==
16
)
?
32
'h
0000ffff
:
(
NUMIRQSRC
==
15
)
?
32
'h
00007fff
:
(
NUMIRQSRC
==
14
)
?
32
'h
00003fff
:
(
NUMIRQSRC
==
13
)
?
32
'h
00001fff
:
(
NUMIRQSRC
==
12
)
?
32
'h
00000fff
:
(
NUMIRQSRC
==
11
)
?
32
'h
000007ff
:
(
NUMIRQSRC
==
10
)
?
32
'h
000003ff
:
(
NUMIRQSRC
==
9
)
?
32
'h
000001ff
:
(
NUMIRQSRC
==
8
)
?
32
'h
000000ff
:
(
NUMIRQSRC
==
7
)
?
32
'h
0000007f
:
(
NUMIRQSRC
==
6
)
?
32
'h
0000003f
:
(
NUMIRQSRC
==
5
)
?
32
'h
0000001f
:
(
NUMIRQSRC
==
4
)
?
32
'h
0000000f
:
(
NUMIRQSRC
==
3
)
?
32
'h
00000007
:
(
NUMIRQSRC
==
2
)
?
32
'h
00000003
:
(
NUMIRQSRC
==
1
)
?
32
'h
00000001
:
(
NUMIRQSRC
==
0
)
?
32
'h
00000000
:
32
'h
00000000
;
assign
CoreInterrupt_l0I
=
CoreInterrupt_I1
&
CoreInterrupt_III
;
assign
CoreInterrupt_lOl
=
PWDATA
&
CoreInterrupt_III
;
assign
CoreInterrupt_OII
=
(
NUMFIQSRC
==
8
)
?
8
'h
ff
:
(
NUMFIQSRC
==
7
)
?
8
'h
7f
:
(
NUMFIQSRC
==
6
)
?
8
'h
3f
:
(
NUMFIQSRC
==
5
)
?
8
'h
1f
:
(
NUMFIQSRC
==
4
)
?
8
'h
0f
:
(
NUMFIQSRC
==
3
)
?
8
'h
07
:
(
NUMFIQSRC
==
2
)
?
8
'h
03
:
(
NUMFIQSRC
==
1
)
?
8
'h
01
:
(
NUMFIQSRC
==
0
)
?
8
'h
00
:
8
'h
00
;
assign
CoreInterrupt_OlI
=
CoreInterrupt_O1
&
CoreInterrupt_OII
;
assign
CoreInterrupt_IOl
=
PWDATA
[
7
:
0
]
&
CoreInterrupt_OII
;
assign
CoreInterrupt_IlI
=
CoreInterrupt_OlI
|
CoreInterrupt_O0I
;
assign
CoreInterrupt_llI
=
CoreInterrupt_IlI
&
CoreInterrupt_I0I
;
assign
FIQ
=
(
FIQPOLARITY
==
1
)
?
|
(
CoreInterrupt_llI
)
:
!
(
|
(
CoreInterrupt_llI
)
)
;
assign
CoreInterrupt_O1I
=
CoreInterrupt_l0I
|
CoreInterrupt_l1I
;
assign
CoreInterrupt_I1I
=
CoreInterrupt_O1I
&
CoreInterrupt_OOl
;
assign
IRQ
=
(
IRQPOLARITY
==
1
)
?
|
(
CoreInterrupt_I1I
)
:
!
(
|
(
CoreInterrupt_I1I
)
)
;
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
if
(
!
PRESETn
)
CoreInterrupt_O0I
<=
{
8
{
1
'b
0
}
}
;
else
if
(
CoreInterrupt_lII
)
case
(
PADDR
)
`CoreInterrupt_O
:
CoreInterrupt_O0I
<=
(
CoreInterrupt_O0I
|
CoreInterrupt_IOl
)
;
`CoreInterrupt_I
:
CoreInterrupt_O0I
<=
(
CoreInterrupt_O0I
&
~
CoreInterrupt_IOl
)
;
default
:
CoreInterrupt_O0I
<=
CoreInterrupt_O0I
;
endcase
end
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
if
(
!
PRESETn
)
CoreInterrupt_I0I
<=
{
8
{
1
'b
0
}
}
;
else
if
(
CoreInterrupt_lII
)
case
(
PADDR
)
`CoreInterrupt_l
:
CoreInterrupt_I0I
<=
(
CoreInterrupt_I0I
|
CoreInterrupt_IOl
)
;
`CoreInterrupt_OI
:
CoreInterrupt_I0I
<=
(
CoreInterrupt_I0I
&
~
CoreInterrupt_IOl
)
;
default
:
CoreInterrupt_I0I
<=
CoreInterrupt_I0I
;
endcase
end
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
if
(
!
PRESETn
)
CoreInterrupt_l1I
<=
{
32
{
1
'b
0
}
}
;
else
if
(
CoreInterrupt_lII
)
case
(
PADDR
)
`CoreInterrupt_Ol
:
CoreInterrupt_l1I
<=
(
CoreInterrupt_l1I
|
CoreInterrupt_lOl
)
;
`CoreInterrupt_Il
:
CoreInterrupt_l1I
<=
(
CoreInterrupt_l1I
&
~
CoreInterrupt_lOl
)
;
default
:
CoreInterrupt_l1I
<=
CoreInterrupt_l1I
;
endcase
end
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
if
(
!
PRESETn
)
CoreInterrupt_OOl
<=
{
32
{
1
'b
0
}
}
;
else
if
(
CoreInterrupt_lII
)
case
(
PADDR
)
`CoreInterrupt_ll
:
CoreInterrupt_OOl
<=
(
CoreInterrupt_OOl
|
CoreInterrupt_lOl
)
;
`CoreInterrupt_O0
:
CoreInterrupt_OOl
<=
(
CoreInterrupt_OOl
&
~
CoreInterrupt_lOl
)
;
default
:
CoreInterrupt_OOl
<=
CoreInterrupt_OOl
;
endcase
end
always
@
(
PSEL
or
PWRITE
or
PADDR
or
CoreInterrupt_O0I
or
CoreInterrupt_I0I
or
CoreInterrupt_IlI
or
CoreInterrupt_llI
or
CoreInterrupt_l1I
or
CoreInterrupt_OOl
or
CoreInterrupt_O1I
or
CoreInterrupt_I1I
)
begin
:
CoreInterrupt_OIl
CoreInterrupt_lOI
=
{
32
{
1
'b
0
}
}
;
if
(
!
PWRITE
&&
PSEL
)
case
(
PADDR
)
`CoreInterrupt_O
:
CoreInterrupt_lOI
[
7
:
0
]
=
CoreInterrupt_O0I
;
`CoreInterrupt_l
:
CoreInterrupt_lOI
[
7
:
0
]
=
CoreInterrupt_I0I
;
`CoreInterrupt_II
:
CoreInterrupt_lOI
[
7
:
0
]
=
CoreInterrupt_IlI
;
`CoreInterrupt_lI
:
CoreInterrupt_lOI
[
7
:
0
]
=
CoreInterrupt_llI
;
`CoreInterrupt_Ol
:
CoreInterrupt_lOI
[
31
:
0
]
=
CoreInterrupt_l1I
;
`CoreInterrupt_ll
:
CoreInterrupt_lOI
[
31
:
0
]
=
CoreInterrupt_OOl
;
`CoreInterrupt_I0
:
CoreInterrupt_lOI
[
31
:
0
]
=
CoreInterrupt_O1I
;
`CoreInterrupt_l0
:
CoreInterrupt_lOI
[
31
:
0
]
=
CoreInterrupt_I1I
;
default
:
CoreInterrupt_lOI
[
31
:
0
]
=
{
32
{
1
'b
0
}
}
;
endcase
else
CoreInterrupt_lOI
=
{
32
{
1
'b
0
}
}
;
end
assign
CoreInterrupt_IOI
=
(
PSEL
&&
!
PWRITE
&&
!
PENABLE
)
;
assign
CoreInterrupt_l1
=
(
CoreInterrupt_IOI
)
?
CoreInterrupt_lOI
:
{
32
{
1
'b
0
}
}
;
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreInterrupt_IIl
if
(
!
PRESETn
)
CoreInterrupt_OOI
<=
{
32
{
1
'b
0
}
}
;
else
CoreInterrupt_OOI
<=
CoreInterrupt_l1
;
end
assign
PRDATA
=
CoreInterrupt_OOI
;
endmodule
