library verilog;
use verilog.vl_types.all;
entity BFM_MAIN is
    generic(
        OPMODE          : integer := 0;
        VECTFILE        : string  := "test.vec";
        MAX_INSTRUCTIONS: integer := 16384;
        MAX_STACK       : integer := 1024;
        MAX_MEMTEST     : integer := 65536;
        TPD             : integer := 1;
        DEBUGLEVEL      : integer := -1;
        CON_SPULSE      : integer := 0;
        ARGVALUE0       : integer := 0;
        ARGVALUE1       : integer := 0;
        ARGVALUE2       : integer := 0;
        ARGVALUE3       : integer := 0;
        ARGVALUE4       : integer := 0;
        ARGVALUE5       : integer := 0;
        ARGVALUE6       : integer := 0;
        ARGVALUE7       : integer := 0;
        ARGVALUE8       : integer := 0;
        ARGVALUE9       : integer := 0;
        ARGVALUE10      : integer := 0;
        ARGVALUE11      : integer := 0;
        ARGVALUE12      : integer := 0;
        ARGVALUE13      : integer := 0;
        ARGVALUE14      : integer := 0;
        ARGVALUE15      : integer := 0;
        ARGVALUE16      : integer := 0;
        ARGVALUE17      : integer := 0;
        ARGVALUE18      : integer := 0;
        ARGVALUE19      : integer := 0;
        ARGVALUE20      : integer := 0;
        ARGVALUE21      : integer := 0;
        ARGVALUE22      : integer := 0;
        ARGVALUE23      : integer := 0;
        ARGVALUE24      : integer := 0;
        ARGVALUE25      : integer := 0;
        ARGVALUE26      : integer := 0;
        ARGVALUE27      : integer := 0;
        ARGVALUE28      : integer := 0;
        ARGVALUE29      : integer := 0;
        ARGVALUE30      : integer := 0;
        ARGVALUE31      : integer := 0;
        ARGVALUE32      : integer := 0;
        ARGVALUE33      : integer := 0;
        ARGVALUE34      : integer := 0;
        ARGVALUE35      : integer := 0;
        ARGVALUE36      : integer := 0;
        ARGVALUE37      : integer := 0;
        ARGVALUE38      : integer := 0;
        ARGVALUE39      : integer := 0;
        ARGVALUE40      : integer := 0;
        ARGVALUE41      : integer := 0;
        ARGVALUE42      : integer := 0;
        ARGVALUE43      : integer := 0;
        ARGVALUE44      : integer := 0;
        ARGVALUE45      : integer := 0;
        ARGVALUE46      : integer := 0;
        ARGVALUE47      : integer := 0;
        ARGVALUE48      : integer := 0;
        ARGVALUE49      : integer := 0;
        ARGVALUE50      : integer := 0;
        ARGVALUE51      : integer := 0;
        ARGVALUE52      : integer := 0;
        ARGVALUE53      : integer := 0;
        ARGVALUE54      : integer := 0;
        ARGVALUE55      : integer := 0;
        ARGVALUE56      : integer := 0;
        ARGVALUE57      : integer := 0;
        ARGVALUE58      : integer := 0;
        ARGVALUE59      : integer := 0;
        ARGVALUE60      : integer := 0;
        ARGVALUE61      : integer := 0;
        ARGVALUE62      : integer := 0;
        ARGVALUE63      : integer := 0;
        ARGVALUE64      : integer := 0;
        ARGVALUE65      : integer := 0;
        ARGVALUE66      : integer := 0;
        ARGVALUE67      : integer := 0;
        ARGVALUE68      : integer := 0;
        ARGVALUE69      : integer := 0;
        ARGVALUE70      : integer := 0;
        ARGVALUE71      : integer := 0;
        ARGVALUE72      : integer := 0;
        ARGVALUE73      : integer := 0;
        ARGVALUE74      : integer := 0;
        ARGVALUE75      : integer := 0;
        ARGVALUE76      : integer := 0;
        ARGVALUE77      : integer := 0;
        ARGVALUE78      : integer := 0;
        ARGVALUE79      : integer := 0;
        ARGVALUE80      : integer := 0;
        ARGVALUE81      : integer := 0;
        ARGVALUE82      : integer := 0;
        ARGVALUE83      : integer := 0;
        ARGVALUE84      : integer := 0;
        ARGVALUE85      : integer := 0;
        ARGVALUE86      : integer := 0;
        ARGVALUE87      : integer := 0;
        ARGVALUE88      : integer := 0;
        ARGVALUE89      : integer := 0;
        ARGVALUE90      : integer := 0;
        ARGVALUE91      : integer := 0;
        ARGVALUE92      : integer := 0;
        ARGVALUE93      : integer := 0;
        ARGVALUE94      : integer := 0;
        ARGVALUE95      : integer := 0;
        ARGVALUE96      : integer := 0;
        ARGVALUE97      : integer := 0;
        ARGVALUE98      : integer := 0;
        ARGVALUE99      : integer := 0;
        ZEROLV          : integer := 0;
        ZERO256         : integer := 0;
        idle            : integer := 0;
        init            : integer := 1;
        active          : integer := 2;
        done            : integer := 3;
        fill            : integer := 4;
        scan            : integer := 5
    );
    port(
        SYSCLK          : in     vl_logic;
        SYSRSTN         : in     vl_logic;
        PCLK            : out    vl_logic;
        HCLK            : out    vl_logic;
        HRESETN         : out    vl_logic;
        HADDR           : out    vl_logic_vector(31 downto 0);
        HBURST          : out    vl_logic_vector(2 downto 0);
        HMASTLOCK       : out    vl_logic;
        HPROT           : out    vl_logic_vector(3 downto 0);
        HSIZE           : out    vl_logic_vector(2 downto 0);
        HTRANS          : out    vl_logic_vector(1 downto 0);
        HWRITE          : out    vl_logic;
        HWDATA          : out    vl_logic_vector(31 downto 0);
        HRDATA          : in     vl_logic_vector(31 downto 0);
        HREADY          : in     vl_logic;
        HRESP           : in     vl_logic;
        HSEL            : out    vl_logic_vector(15 downto 0);
        INTERRUPT       : in     vl_logic_vector(255 downto 0);
        GP_OUT          : out    vl_logic_vector(31 downto 0);
        GP_IN           : in     vl_logic_vector(31 downto 0);
        EXT_WR          : out    vl_logic;
        EXT_RD          : out    vl_logic;
        EXT_ADDR        : out    vl_logic_vector(31 downto 0);
        EXT_DATA        : inout  vl_logic_vector(31 downto 0);
        EXT_WAIT        : in     vl_logic;
        CON_ADDR        : in     vl_logic_vector(15 downto 0);
        CON_DATA        : inout  vl_logic_vector(31 downto 0);
        CON_RD          : in     vl_logic;
        CON_WR          : in     vl_logic;
        CON_BUSY        : out    vl_logic;
        INSTR_OUT       : out    vl_logic_vector(31 downto 0);
        INSTR_IN        : in     vl_logic_vector(31 downto 0);
        FINISHED        : out    vl_logic;
        FAILED          : out    vl_logic
    );
end BFM_MAIN;
