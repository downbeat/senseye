library verilog;
use verilog.vl_types.all;
entity F2DSS_SSE_ENGINE is
    generic(
        RAM_DEBUG       : integer := 0
    );
    port(
        PRESETN         : in     vl_logic;
        PCLK            : in     vl_logic;
        TDM_CNT         : in     vl_logic_vector(2 downto 0);
        SSE_TS_CTRL0    : out    vl_logic;
        SSE_RWB         : in     vl_logic;
        SSE_ADDR        : in     vl_logic_vector(9 downto 0);
        SSE_WDATA       : in     vl_logic_vector(15 downto 0);
        SSE_RDATA_o     : out    vl_logic_vector(15 downto 0);
        PPE_FIFO_FULL   : in     vl_logic;
        PC0_FLAGS_o     : out    vl_logic_vector(3 downto 0);
        PC1_FLAGS_o     : out    vl_logic_vector(3 downto 0);
        PC2_FLAGS_o     : out    vl_logic_vector(3 downto 0);
        ADC0_CALIBRATE_rise: out    vl_logic;
        ADC1_CALIBRATE_rise: out    vl_logic;
        ADC2_CALIBRATE_rise: out    vl_logic;
        ADC0_CALIBRATE_fall: out    vl_logic;
        ADC1_CALIBRATE_fall: out    vl_logic;
        ADC2_CALIBRATE_fall: out    vl_logic;
        ADC0_DATAVALID_rise: out    vl_logic;
        ADC1_DATAVALID_rise: out    vl_logic;
        ADC2_DATAVALID_rise: out    vl_logic;
        ADC0_BUSY       : in     vl_logic;
        ADC1_BUSY       : in     vl_logic;
        ADC2_BUSY       : in     vl_logic;
        ADC0_CALIBRATE  : in     vl_logic;
        ADC1_CALIBRATE  : in     vl_logic;
        ADC2_CALIBRATE  : in     vl_logic;
        ADC0_DATAVALID  : in     vl_logic;
        ADC1_DATAVALID  : in     vl_logic;
        ADC2_DATAVALID  : in     vl_logic;
        ADC0_SAMPLE     : in     vl_logic;
        ADC1_SAMPLE     : in     vl_logic;
        ADC2_SAMPLE     : in     vl_logic;
        ADC0_TVC_o      : out    vl_logic_vector(7 downto 0);
        ADC1_TVC_o      : out    vl_logic_vector(7 downto 0);
        ADC2_TVC_o      : out    vl_logic_vector(7 downto 0);
        ADC0_STC_o      : out    vl_logic_vector(7 downto 0);
        ADC1_STC_o      : out    vl_logic_vector(7 downto 0);
        ADC2_STC_o      : out    vl_logic_vector(7 downto 0);
        ADC0_MODE_o     : out    vl_logic_vector(3 downto 0);
        ADC1_MODE_o     : out    vl_logic_vector(3 downto 0);
        ADC2_MODE_o     : out    vl_logic_vector(3 downto 0);
        ADC_VAREFSEL_o  : out    vl_logic;
        ABPOWERON_o     : out    vl_logic;
        ADC0_CHNUMBER_o : out    vl_logic_vector(4 downto 0);
        ADC1_CHNUMBER_o : out    vl_logic_vector(4 downto 0);
        ADC2_CHNUMBER_o : out    vl_logic_vector(4 downto 0);
        ADC0_ADCSTART_o : out    vl_logic;
        ADC1_ADCSTART_o : out    vl_logic;
        ADC2_ADCSTART_o : out    vl_logic;
        ADC0_PWRDWN_o   : out    vl_logic;
        ADC1_PWRDWN_o   : out    vl_logic;
        ADC2_PWRDWN_o   : out    vl_logic;
        ADC0_ADCRESET_o : out    vl_logic;
        ADC1_ADCRESET_o : out    vl_logic;
        ADC2_ADCRESET_o : out    vl_logic;
        ACB_RDATA       : in     vl_logic_vector(7 downto 0);
        ACB_ADDR        : out    vl_logic_vector(7 downto 0);
        ACB_WRE         : out    vl_logic;
        ACB_WDATA       : out    vl_logic_vector(7 downto 0);
        ACB_RESETN      : out    vl_logic;
        DAC0_DATA_o     : out    vl_logic_vector(23 downto 0);
        DAC1_DATA_o     : out    vl_logic_vector(23 downto 0);
        DAC2_DATA_o     : out    vl_logic_vector(23 downto 0);
        DAC0_CTRL_o     : out    vl_logic_vector(7 downto 0);
        DAC1_CTRL_o     : out    vl_logic_vector(7 downto 0);
        DAC2_CTRL_o     : out    vl_logic_vector(7 downto 0);
        PDMA_decode     : in     vl_logic;
        INREADY_o       : out    vl_logic;
        SSE_ADC0_RESULTS_o: out    vl_logic;
        SSE_ADC1_RESULTS_o: out    vl_logic;
        SSE_ADC2_RESULTS_o: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of RAM_DEBUG : constant is 1;
end F2DSS_SSE_ENGINE;
